// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 18 2025 11:07:06

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    generated_signal,
    RST_N,
    ENdin,
    CLK);

    output generated_signal;
    input RST_N;
    output ENdin;
    input CLK;

    wire N__1640;
    wire N__1639;
    wire N__1638;
    wire N__1629;
    wire N__1628;
    wire N__1627;
    wire N__1620;
    wire N__1619;
    wire N__1618;
    wire N__1611;
    wire N__1610;
    wire N__1609;
    wire N__1592;
    wire N__1589;
    wire N__1588;
    wire N__1587;
    wire N__1584;
    wire N__1581;
    wire N__1578;
    wire N__1571;
    wire N__1568;
    wire N__1565;
    wire N__1564;
    wire N__1563;
    wire N__1558;
    wire N__1555;
    wire N__1550;
    wire N__1547;
    wire N__1546;
    wire N__1543;
    wire N__1540;
    wire N__1535;
    wire N__1532;
    wire N__1531;
    wire N__1530;
    wire N__1527;
    wire N__1522;
    wire N__1519;
    wire N__1514;
    wire N__1511;
    wire N__1510;
    wire N__1507;
    wire N__1504;
    wire N__1499;
    wire N__1496;
    wire N__1495;
    wire N__1492;
    wire N__1489;
    wire N__1486;
    wire N__1481;
    wire N__1478;
    wire N__1477;
    wire N__1476;
    wire N__1475;
    wire N__1474;
    wire N__1473;
    wire N__1472;
    wire N__1471;
    wire N__1462;
    wire N__1453;
    wire N__1448;
    wire N__1445;
    wire N__1444;
    wire N__1441;
    wire N__1438;
    wire N__1433;
    wire N__1432;
    wire N__1431;
    wire N__1430;
    wire N__1429;
    wire N__1428;
    wire N__1427;
    wire N__1426;
    wire N__1425;
    wire N__1424;
    wire N__1423;
    wire N__1422;
    wire N__1397;
    wire N__1394;
    wire N__1391;
    wire N__1390;
    wire N__1389;
    wire N__1388;
    wire N__1387;
    wire N__1386;
    wire N__1385;
    wire N__1384;
    wire N__1367;
    wire N__1364;
    wire N__1361;
    wire N__1358;
    wire N__1355;
    wire N__1352;
    wire N__1349;
    wire N__1346;
    wire N__1343;
    wire N__1340;
    wire N__1337;
    wire N__1334;
    wire N__1331;
    wire N__1328;
    wire N__1325;
    wire N__1322;
    wire N__1319;
    wire N__1318;
    wire N__1317;
    wire N__1316;
    wire N__1315;
    wire N__1314;
    wire N__1313;
    wire N__1310;
    wire N__1297;
    wire N__1296;
    wire N__1295;
    wire N__1294;
    wire N__1293;
    wire N__1292;
    wire N__1291;
    wire N__1290;
    wire N__1289;
    wire N__1286;
    wire N__1283;
    wire N__1266;
    wire N__1259;
    wire N__1256;
    wire N__1253;
    wire N__1250;
    wire N__1247;
    wire N__1246;
    wire N__1243;
    wire N__1240;
    wire N__1235;
    wire N__1234;
    wire N__1233;
    wire N__1228;
    wire N__1225;
    wire N__1220;
    wire N__1217;
    wire N__1216;
    wire N__1211;
    wire N__1208;
    wire N__1207;
    wire N__1206;
    wire N__1205;
    wire N__1202;
    wire N__1199;
    wire N__1194;
    wire N__1187;
    wire N__1186;
    wire N__1183;
    wire N__1180;
    wire N__1175;
    wire N__1172;
    wire N__1169;
    wire N__1166;
    wire N__1163;
    wire N__1160;
    wire N__1157;
    wire N__1154;
    wire N__1151;
    wire N__1148;
    wire N__1145;
    wire N__1142;
    wire N__1139;
    wire N__1136;
    wire N__1133;
    wire N__1130;
    wire N__1127;
    wire N__1124;
    wire N__1121;
    wire N__1118;
    wire N__1115;
    wire N__1112;
    wire N__1109;
    wire N__1108;
    wire N__1107;
    wire N__1106;
    wire N__1097;
    wire N__1094;
    wire N__1093;
    wire N__1092;
    wire N__1091;
    wire N__1090;
    wire N__1089;
    wire N__1086;
    wire N__1083;
    wire N__1072;
    wire N__1067;
    wire N__1066;
    wire N__1065;
    wire N__1064;
    wire N__1061;
    wire N__1060;
    wire N__1049;
    wire N__1046;
    wire N__1045;
    wire N__1044;
    wire N__1043;
    wire N__1040;
    wire N__1039;
    wire N__1036;
    wire N__1035;
    wire N__1034;
    wire N__1033;
    wire N__1032;
    wire N__1029;
    wire N__1026;
    wire N__1023;
    wire N__1010;
    wire N__1001;
    wire N__1000;
    wire N__997;
    wire N__994;
    wire N__993;
    wire N__990;
    wire N__985;
    wire N__982;
    wire N__979;
    wire N__976;
    wire N__973;
    wire N__970;
    wire N__967;
    wire N__964;
    wire N__961;
    wire N__956;
    wire N__955;
    wire N__954;
    wire N__953;
    wire N__952;
    wire N__947;
    wire N__946;
    wire N__945;
    wire N__942;
    wire N__937;
    wire N__934;
    wire N__929;
    wire N__920;
    wire N__919;
    wire N__918;
    wire N__917;
    wire N__914;
    wire N__909;
    wire N__906;
    wire N__899;
    wire N__896;
    wire N__893;
    wire N__892;
    wire N__889;
    wire N__886;
    wire N__881;
    wire N__878;
    wire N__875;
    wire N__872;
    wire N__869;
    wire N__866;
    wire N__863;
    wire N__860;
    wire N__857;
    wire N__854;
    wire N__851;
    wire N__848;
    wire N__845;
    wire N__842;
    wire N__841;
    wire N__838;
    wire N__835;
    wire N__830;
    wire N__827;
    wire N__826;
    wire N__825;
    wire N__822;
    wire N__817;
    wire N__814;
    wire N__809;
    wire N__806;
    wire N__803;
    wire N__800;
    wire N__799;
    wire N__798;
    wire N__797;
    wire N__796;
    wire N__791;
    wire N__784;
    wire N__779;
    wire N__778;
    wire N__777;
    wire N__776;
    wire N__769;
    wire N__766;
    wire N__763;
    wire N__758;
    wire N__755;
    wire N__754;
    wire N__753;
    wire N__750;
    wire N__749;
    wire N__746;
    wire N__743;
    wire N__742;
    wire N__737;
    wire N__730;
    wire N__725;
    wire N__722;
    wire N__719;
    wire N__716;
    wire VCCG0;
    wire GNDG0;
    wire RST_N_c_i;
    wire \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_ ;
    wire \fsm_shiftRegs_inst1.counterZ0Z_0 ;
    wire \fsm_shiftRegs_inst1.counterZ0Z_1 ;
    wire \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3_cascade_ ;
    wire \fsm_shiftRegs_inst1.counterZ0Z_3 ;
    wire ENdin_c;
    wire enable_din;
    wire \fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_ ;
    wire \fsm_shiftRegs_inst1.N_123_1 ;
    wire \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_ ;
    wire \fsm_shiftRegs_inst1.counterDYNZ0Z_3 ;
    wire \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3 ;
    wire \fsm_shiftRegs_inst1.counterDYNZ0Z_2 ;
    wire \fsm_shiftRegs_inst1.counterDYNZ0Z_0 ;
    wire \fsm_shiftRegs_inst1.counterDYNZ0Z_1 ;
    wire \fsm_shiftRegs_inst1.current_stateZ0Z_2 ;
    wire RST_N_c;
    wire \fsm_shiftRegs_inst1.current_stateZ0Z_1 ;
    wire \fsm_shiftRegs_inst1.counterZ0Z_2 ;
    wire \fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2 ;
    wire \fsm_shiftRegs_inst1.current_stateZ0Z_3 ;
    wire \fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_ ;
    wire \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_ ;
    wire \fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0 ;
    wire \fsm_shiftRegs_inst1.current_stateZ0Z_4 ;
    wire signal_out_fsm;
    wire SELSTAT;
    wire SELDYN;
    wire generated_signal_c;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_2 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_3 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_6 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_4 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_5 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_15 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_11 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_12 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_10 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_13 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_14 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_9 ;
    wire \fsm_shiftRegs_inst1.current_stateZ0Z_0 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_7 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_8 ;
    wire \fsm_shiftRegs_inst1.un1_current_state4_0 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_0 ;
    wire bfn_14_15_0_;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_1 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_0 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_2 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_1 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_3 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_2 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_4 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_3 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_5 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_4 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_6 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_5 ;
    wire \fsm_shiftRegs_inst1.current_state_i_4 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_6 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_7 ;
    wire _gnd_net_;
    wire CLK_c_g;
    wire RST_N_c_i_g;

    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__1638),
            .GLOBALBUFFEROUTPUT(CLK_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__1640),
            .DIN(N__1639),
            .DOUT(N__1638),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__1640),
            .PADOUT(N__1639),
            .PADIN(N__1638),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RST_N_ibuf_iopad (
            .OE(N__1629),
            .DIN(N__1628),
            .DOUT(N__1627),
            .PACKAGEPIN(RST_N));
    defparam RST_N_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RST_N_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RST_N_ibuf_preio (
            .PADOEN(N__1629),
            .PADOUT(N__1628),
            .PADIN(N__1627),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RST_N_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD generated_signal_obuf_iopad (
            .OE(N__1620),
            .DIN(N__1619),
            .DOUT(N__1618),
            .PACKAGEPIN(generated_signal));
    defparam generated_signal_obuf_preio.NEG_TRIGGER=1'b0;
    defparam generated_signal_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO generated_signal_obuf_preio (
            .PADOEN(N__1620),
            .PADOUT(N__1619),
            .PADIN(N__1618),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1163),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ENdin_obuf_iopad (
            .OE(N__1611),
            .DIN(N__1610),
            .DOUT(N__1609),
            .PACKAGEPIN(ENdin));
    defparam ENdin_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ENdin_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ENdin_obuf_preio (
            .PADOEN(N__1611),
            .PADOUT(N__1610),
            .PADIN(N__1609),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__875),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__355 (
            .O(N__1592),
            .I(N__1589));
    LocalMux I__354 (
            .O(N__1589),
            .I(N__1584));
    InMux I__353 (
            .O(N__1588),
            .I(N__1581));
    InMux I__352 (
            .O(N__1587),
            .I(N__1578));
    Odrv4 I__351 (
            .O(N__1584),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_1 ));
    LocalMux I__350 (
            .O(N__1581),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_1 ));
    LocalMux I__349 (
            .O(N__1578),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_1 ));
    InMux I__348 (
            .O(N__1571),
            .I(\fsm_shiftRegs_inst1.counter2_cry_0 ));
    CascadeMux I__347 (
            .O(N__1568),
            .I(N__1565));
    InMux I__346 (
            .O(N__1565),
            .I(N__1558));
    InMux I__345 (
            .O(N__1564),
            .I(N__1558));
    InMux I__344 (
            .O(N__1563),
            .I(N__1555));
    LocalMux I__343 (
            .O(N__1558),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_2 ));
    LocalMux I__342 (
            .O(N__1555),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_2 ));
    InMux I__341 (
            .O(N__1550),
            .I(\fsm_shiftRegs_inst1.counter2_cry_1 ));
    InMux I__340 (
            .O(N__1547),
            .I(N__1543));
    InMux I__339 (
            .O(N__1546),
            .I(N__1540));
    LocalMux I__338 (
            .O(N__1543),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_3 ));
    LocalMux I__337 (
            .O(N__1540),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_3 ));
    InMux I__336 (
            .O(N__1535),
            .I(\fsm_shiftRegs_inst1.counter2_cry_2 ));
    CascadeMux I__335 (
            .O(N__1532),
            .I(N__1527));
    InMux I__334 (
            .O(N__1531),
            .I(N__1522));
    InMux I__333 (
            .O(N__1530),
            .I(N__1522));
    InMux I__332 (
            .O(N__1527),
            .I(N__1519));
    LocalMux I__331 (
            .O(N__1522),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_4 ));
    LocalMux I__330 (
            .O(N__1519),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_4 ));
    InMux I__329 (
            .O(N__1514),
            .I(\fsm_shiftRegs_inst1.counter2_cry_3 ));
    InMux I__328 (
            .O(N__1511),
            .I(N__1507));
    InMux I__327 (
            .O(N__1510),
            .I(N__1504));
    LocalMux I__326 (
            .O(N__1507),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_5 ));
    LocalMux I__325 (
            .O(N__1504),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_5 ));
    InMux I__324 (
            .O(N__1499),
            .I(\fsm_shiftRegs_inst1.counter2_cry_4 ));
    CascadeMux I__323 (
            .O(N__1496),
            .I(N__1492));
    InMux I__322 (
            .O(N__1495),
            .I(N__1489));
    InMux I__321 (
            .O(N__1492),
            .I(N__1486));
    LocalMux I__320 (
            .O(N__1489),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_6 ));
    LocalMux I__319 (
            .O(N__1486),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_6 ));
    InMux I__318 (
            .O(N__1481),
            .I(\fsm_shiftRegs_inst1.counter2_cry_5 ));
    InMux I__317 (
            .O(N__1478),
            .I(N__1462));
    InMux I__316 (
            .O(N__1477),
            .I(N__1462));
    InMux I__315 (
            .O(N__1476),
            .I(N__1462));
    InMux I__314 (
            .O(N__1475),
            .I(N__1462));
    InMux I__313 (
            .O(N__1474),
            .I(N__1453));
    InMux I__312 (
            .O(N__1473),
            .I(N__1453));
    InMux I__311 (
            .O(N__1472),
            .I(N__1453));
    InMux I__310 (
            .O(N__1471),
            .I(N__1453));
    LocalMux I__309 (
            .O(N__1462),
            .I(\fsm_shiftRegs_inst1.current_state_i_4 ));
    LocalMux I__308 (
            .O(N__1453),
            .I(\fsm_shiftRegs_inst1.current_state_i_4 ));
    InMux I__307 (
            .O(N__1448),
            .I(\fsm_shiftRegs_inst1.counter2_cry_6 ));
    InMux I__306 (
            .O(N__1445),
            .I(N__1441));
    InMux I__305 (
            .O(N__1444),
            .I(N__1438));
    LocalMux I__304 (
            .O(N__1441),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_7 ));
    LocalMux I__303 (
            .O(N__1438),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_7 ));
    ClkMux I__302 (
            .O(N__1433),
            .I(N__1397));
    ClkMux I__301 (
            .O(N__1432),
            .I(N__1397));
    ClkMux I__300 (
            .O(N__1431),
            .I(N__1397));
    ClkMux I__299 (
            .O(N__1430),
            .I(N__1397));
    ClkMux I__298 (
            .O(N__1429),
            .I(N__1397));
    ClkMux I__297 (
            .O(N__1428),
            .I(N__1397));
    ClkMux I__296 (
            .O(N__1427),
            .I(N__1397));
    ClkMux I__295 (
            .O(N__1426),
            .I(N__1397));
    ClkMux I__294 (
            .O(N__1425),
            .I(N__1397));
    ClkMux I__293 (
            .O(N__1424),
            .I(N__1397));
    ClkMux I__292 (
            .O(N__1423),
            .I(N__1397));
    ClkMux I__291 (
            .O(N__1422),
            .I(N__1397));
    GlobalMux I__290 (
            .O(N__1397),
            .I(N__1394));
    gio2CtrlBuf I__289 (
            .O(N__1394),
            .I(CLK_c_g));
    SRMux I__288 (
            .O(N__1391),
            .I(N__1367));
    SRMux I__287 (
            .O(N__1390),
            .I(N__1367));
    SRMux I__286 (
            .O(N__1389),
            .I(N__1367));
    SRMux I__285 (
            .O(N__1388),
            .I(N__1367));
    SRMux I__284 (
            .O(N__1387),
            .I(N__1367));
    SRMux I__283 (
            .O(N__1386),
            .I(N__1367));
    SRMux I__282 (
            .O(N__1385),
            .I(N__1367));
    SRMux I__281 (
            .O(N__1384),
            .I(N__1367));
    GlobalMux I__280 (
            .O(N__1367),
            .I(N__1364));
    gio2CtrlBuf I__279 (
            .O(N__1364),
            .I(RST_N_c_i_g));
    InMux I__278 (
            .O(N__1361),
            .I(N__1358));
    LocalMux I__277 (
            .O(N__1358),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_15 ));
    InMux I__276 (
            .O(N__1355),
            .I(N__1352));
    LocalMux I__275 (
            .O(N__1352),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_11 ));
    InMux I__274 (
            .O(N__1349),
            .I(N__1346));
    LocalMux I__273 (
            .O(N__1346),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_12 ));
    InMux I__272 (
            .O(N__1343),
            .I(N__1340));
    LocalMux I__271 (
            .O(N__1340),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_10 ));
    InMux I__270 (
            .O(N__1337),
            .I(N__1334));
    LocalMux I__269 (
            .O(N__1334),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_13 ));
    InMux I__268 (
            .O(N__1331),
            .I(N__1328));
    LocalMux I__267 (
            .O(N__1328),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_14 ));
    InMux I__266 (
            .O(N__1325),
            .I(N__1322));
    LocalMux I__265 (
            .O(N__1322),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_9 ));
    CascadeMux I__264 (
            .O(N__1319),
            .I(N__1310));
    InMux I__263 (
            .O(N__1318),
            .I(N__1297));
    InMux I__262 (
            .O(N__1317),
            .I(N__1297));
    InMux I__261 (
            .O(N__1316),
            .I(N__1297));
    InMux I__260 (
            .O(N__1315),
            .I(N__1297));
    InMux I__259 (
            .O(N__1314),
            .I(N__1297));
    InMux I__258 (
            .O(N__1313),
            .I(N__1297));
    InMux I__257 (
            .O(N__1310),
            .I(N__1286));
    LocalMux I__256 (
            .O(N__1297),
            .I(N__1283));
    InMux I__255 (
            .O(N__1296),
            .I(N__1266));
    InMux I__254 (
            .O(N__1295),
            .I(N__1266));
    InMux I__253 (
            .O(N__1294),
            .I(N__1266));
    InMux I__252 (
            .O(N__1293),
            .I(N__1266));
    InMux I__251 (
            .O(N__1292),
            .I(N__1266));
    InMux I__250 (
            .O(N__1291),
            .I(N__1266));
    InMux I__249 (
            .O(N__1290),
            .I(N__1266));
    InMux I__248 (
            .O(N__1289),
            .I(N__1266));
    LocalMux I__247 (
            .O(N__1286),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_0 ));
    Odrv4 I__246 (
            .O(N__1283),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_0 ));
    LocalMux I__245 (
            .O(N__1266),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_0 ));
    InMux I__244 (
            .O(N__1259),
            .I(N__1256));
    LocalMux I__243 (
            .O(N__1256),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_7 ));
    InMux I__242 (
            .O(N__1253),
            .I(N__1250));
    LocalMux I__241 (
            .O(N__1250),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_8 ));
    CEMux I__240 (
            .O(N__1247),
            .I(N__1243));
    CEMux I__239 (
            .O(N__1246),
            .I(N__1240));
    LocalMux I__238 (
            .O(N__1243),
            .I(\fsm_shiftRegs_inst1.un1_current_state4_0 ));
    LocalMux I__237 (
            .O(N__1240),
            .I(\fsm_shiftRegs_inst1.un1_current_state4_0 ));
    InMux I__236 (
            .O(N__1235),
            .I(N__1228));
    InMux I__235 (
            .O(N__1234),
            .I(N__1228));
    InMux I__234 (
            .O(N__1233),
            .I(N__1225));
    LocalMux I__233 (
            .O(N__1228),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_0 ));
    LocalMux I__232 (
            .O(N__1225),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_0 ));
    InMux I__231 (
            .O(N__1220),
            .I(bfn_14_15_0_));
    InMux I__230 (
            .O(N__1217),
            .I(N__1211));
    InMux I__229 (
            .O(N__1216),
            .I(N__1211));
    LocalMux I__228 (
            .O(N__1211),
            .I(\fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0 ));
    InMux I__227 (
            .O(N__1208),
            .I(N__1202));
    InMux I__226 (
            .O(N__1207),
            .I(N__1199));
    InMux I__225 (
            .O(N__1206),
            .I(N__1194));
    InMux I__224 (
            .O(N__1205),
            .I(N__1194));
    LocalMux I__223 (
            .O(N__1202),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_4 ));
    LocalMux I__222 (
            .O(N__1199),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_4 ));
    LocalMux I__221 (
            .O(N__1194),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_4 ));
    InMux I__220 (
            .O(N__1187),
            .I(N__1183));
    InMux I__219 (
            .O(N__1186),
            .I(N__1180));
    LocalMux I__218 (
            .O(N__1183),
            .I(signal_out_fsm));
    LocalMux I__217 (
            .O(N__1180),
            .I(signal_out_fsm));
    InMux I__216 (
            .O(N__1175),
            .I(N__1172));
    LocalMux I__215 (
            .O(N__1172),
            .I(SELSTAT));
    InMux I__214 (
            .O(N__1169),
            .I(N__1166));
    LocalMux I__213 (
            .O(N__1166),
            .I(SELDYN));
    IoInMux I__212 (
            .O(N__1163),
            .I(N__1160));
    LocalMux I__211 (
            .O(N__1160),
            .I(N__1157));
    Span4Mux_s1_v I__210 (
            .O(N__1157),
            .I(N__1154));
    Span4Mux_v I__209 (
            .O(N__1154),
            .I(N__1151));
    Sp12to4 I__208 (
            .O(N__1151),
            .I(N__1148));
    Span12Mux_s10_h I__207 (
            .O(N__1148),
            .I(N__1145));
    Span12Mux_v I__206 (
            .O(N__1145),
            .I(N__1142));
    Odrv12 I__205 (
            .O(N__1142),
            .I(generated_signal_c));
    InMux I__204 (
            .O(N__1139),
            .I(N__1136));
    LocalMux I__203 (
            .O(N__1136),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_2 ));
    InMux I__202 (
            .O(N__1133),
            .I(N__1130));
    LocalMux I__201 (
            .O(N__1130),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_3 ));
    InMux I__200 (
            .O(N__1127),
            .I(N__1124));
    LocalMux I__199 (
            .O(N__1124),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_6 ));
    InMux I__198 (
            .O(N__1121),
            .I(N__1118));
    LocalMux I__197 (
            .O(N__1118),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_4 ));
    InMux I__196 (
            .O(N__1115),
            .I(N__1112));
    LocalMux I__195 (
            .O(N__1112),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_5 ));
    InMux I__194 (
            .O(N__1109),
            .I(N__1097));
    InMux I__193 (
            .O(N__1108),
            .I(N__1097));
    InMux I__192 (
            .O(N__1107),
            .I(N__1097));
    InMux I__191 (
            .O(N__1106),
            .I(N__1097));
    LocalMux I__190 (
            .O(N__1097),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_2 ));
    CascadeMux I__189 (
            .O(N__1094),
            .I(N__1086));
    InMux I__188 (
            .O(N__1093),
            .I(N__1083));
    InMux I__187 (
            .O(N__1092),
            .I(N__1072));
    InMux I__186 (
            .O(N__1091),
            .I(N__1072));
    InMux I__185 (
            .O(N__1090),
            .I(N__1072));
    InMux I__184 (
            .O(N__1089),
            .I(N__1072));
    InMux I__183 (
            .O(N__1086),
            .I(N__1072));
    LocalMux I__182 (
            .O(N__1083),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_0 ));
    LocalMux I__181 (
            .O(N__1072),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_0 ));
    CascadeMux I__180 (
            .O(N__1067),
            .I(N__1061));
    InMux I__179 (
            .O(N__1066),
            .I(N__1049));
    InMux I__178 (
            .O(N__1065),
            .I(N__1049));
    InMux I__177 (
            .O(N__1064),
            .I(N__1049));
    InMux I__176 (
            .O(N__1061),
            .I(N__1049));
    InMux I__175 (
            .O(N__1060),
            .I(N__1049));
    LocalMux I__174 (
            .O(N__1049),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_1 ));
    InMux I__173 (
            .O(N__1046),
            .I(N__1040));
    CascadeMux I__172 (
            .O(N__1045),
            .I(N__1036));
    InMux I__171 (
            .O(N__1044),
            .I(N__1029));
    InMux I__170 (
            .O(N__1043),
            .I(N__1026));
    LocalMux I__169 (
            .O(N__1040),
            .I(N__1023));
    InMux I__168 (
            .O(N__1039),
            .I(N__1010));
    InMux I__167 (
            .O(N__1036),
            .I(N__1010));
    InMux I__166 (
            .O(N__1035),
            .I(N__1010));
    InMux I__165 (
            .O(N__1034),
            .I(N__1010));
    InMux I__164 (
            .O(N__1033),
            .I(N__1010));
    InMux I__163 (
            .O(N__1032),
            .I(N__1010));
    LocalMux I__162 (
            .O(N__1029),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ));
    LocalMux I__161 (
            .O(N__1026),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ));
    Odrv4 I__160 (
            .O(N__1023),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ));
    LocalMux I__159 (
            .O(N__1010),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ));
    InMux I__158 (
            .O(N__1001),
            .I(N__997));
    CascadeMux I__157 (
            .O(N__1000),
            .I(N__994));
    LocalMux I__156 (
            .O(N__997),
            .I(N__990));
    InMux I__155 (
            .O(N__994),
            .I(N__985));
    InMux I__154 (
            .O(N__993),
            .I(N__985));
    Sp12to4 I__153 (
            .O(N__990),
            .I(N__982));
    LocalMux I__152 (
            .O(N__985),
            .I(N__979));
    Span12Mux_v I__151 (
            .O(N__982),
            .I(N__976));
    Sp12to4 I__150 (
            .O(N__979),
            .I(N__973));
    Span12Mux_h I__149 (
            .O(N__976),
            .I(N__970));
    Span12Mux_v I__148 (
            .O(N__973),
            .I(N__967));
    Span12Mux_h I__147 (
            .O(N__970),
            .I(N__964));
    Span12Mux_h I__146 (
            .O(N__967),
            .I(N__961));
    Odrv12 I__145 (
            .O(N__964),
            .I(RST_N_c));
    Odrv12 I__144 (
            .O(N__961),
            .I(RST_N_c));
    InMux I__143 (
            .O(N__956),
            .I(N__947));
    InMux I__142 (
            .O(N__955),
            .I(N__947));
    InMux I__141 (
            .O(N__954),
            .I(N__942));
    InMux I__140 (
            .O(N__953),
            .I(N__937));
    InMux I__139 (
            .O(N__952),
            .I(N__937));
    LocalMux I__138 (
            .O(N__947),
            .I(N__934));
    InMux I__137 (
            .O(N__946),
            .I(N__929));
    InMux I__136 (
            .O(N__945),
            .I(N__929));
    LocalMux I__135 (
            .O(N__942),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_1 ));
    LocalMux I__134 (
            .O(N__937),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_1 ));
    Odrv4 I__133 (
            .O(N__934),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_1 ));
    LocalMux I__132 (
            .O(N__929),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_1 ));
    InMux I__131 (
            .O(N__920),
            .I(N__914));
    InMux I__130 (
            .O(N__919),
            .I(N__909));
    InMux I__129 (
            .O(N__918),
            .I(N__909));
    InMux I__128 (
            .O(N__917),
            .I(N__906));
    LocalMux I__127 (
            .O(N__914),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_2 ));
    LocalMux I__126 (
            .O(N__909),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_2 ));
    LocalMux I__125 (
            .O(N__906),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_2 ));
    InMux I__124 (
            .O(N__899),
            .I(N__896));
    LocalMux I__123 (
            .O(N__896),
            .I(\fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2 ));
    InMux I__122 (
            .O(N__893),
            .I(N__889));
    InMux I__121 (
            .O(N__892),
            .I(N__886));
    LocalMux I__120 (
            .O(N__889),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_3 ));
    LocalMux I__119 (
            .O(N__886),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_3 ));
    CascadeMux I__118 (
            .O(N__881),
            .I(\fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_ ));
    CascadeMux I__117 (
            .O(N__878),
            .I(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_ ));
    IoInMux I__116 (
            .O(N__875),
            .I(N__872));
    LocalMux I__115 (
            .O(N__872),
            .I(N__869));
    IoSpan4Mux I__114 (
            .O(N__869),
            .I(N__866));
    Sp12to4 I__113 (
            .O(N__866),
            .I(N__863));
    Span12Mux_s7_h I__112 (
            .O(N__863),
            .I(N__860));
    Span12Mux_h I__111 (
            .O(N__860),
            .I(N__857));
    Odrv12 I__110 (
            .O(N__857),
            .I(ENdin_c));
    InMux I__109 (
            .O(N__854),
            .I(N__851));
    LocalMux I__108 (
            .O(N__851),
            .I(enable_din));
    CascadeMux I__107 (
            .O(N__848),
            .I(\fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_ ));
    InMux I__106 (
            .O(N__845),
            .I(N__842));
    LocalMux I__105 (
            .O(N__842),
            .I(N__838));
    InMux I__104 (
            .O(N__841),
            .I(N__835));
    Odrv4 I__103 (
            .O(N__838),
            .I(\fsm_shiftRegs_inst1.N_123_1 ));
    LocalMux I__102 (
            .O(N__835),
            .I(\fsm_shiftRegs_inst1.N_123_1 ));
    CascadeMux I__101 (
            .O(N__830),
            .I(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_ ));
    CascadeMux I__100 (
            .O(N__827),
            .I(N__822));
    InMux I__99 (
            .O(N__826),
            .I(N__817));
    InMux I__98 (
            .O(N__825),
            .I(N__817));
    InMux I__97 (
            .O(N__822),
            .I(N__814));
    LocalMux I__96 (
            .O(N__817),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_3 ));
    LocalMux I__95 (
            .O(N__814),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_3 ));
    InMux I__94 (
            .O(N__809),
            .I(N__806));
    LocalMux I__93 (
            .O(N__806),
            .I(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3 ));
    CascadeMux I__92 (
            .O(N__803),
            .I(\fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_ ));
    InMux I__91 (
            .O(N__800),
            .I(N__791));
    InMux I__90 (
            .O(N__799),
            .I(N__791));
    InMux I__89 (
            .O(N__798),
            .I(N__784));
    InMux I__88 (
            .O(N__797),
            .I(N__784));
    InMux I__87 (
            .O(N__796),
            .I(N__784));
    LocalMux I__86 (
            .O(N__791),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_0 ));
    LocalMux I__85 (
            .O(N__784),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_0 ));
    InMux I__84 (
            .O(N__779),
            .I(N__769));
    InMux I__83 (
            .O(N__778),
            .I(N__769));
    InMux I__82 (
            .O(N__777),
            .I(N__769));
    InMux I__81 (
            .O(N__776),
            .I(N__766));
    LocalMux I__80 (
            .O(N__769),
            .I(N__763));
    LocalMux I__79 (
            .O(N__766),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_1 ));
    Odrv4 I__78 (
            .O(N__763),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_1 ));
    CascadeMux I__77 (
            .O(N__758),
            .I(\fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3_cascade_ ));
    CascadeMux I__76 (
            .O(N__755),
            .I(N__750));
    CascadeMux I__75 (
            .O(N__754),
            .I(N__746));
    CascadeMux I__74 (
            .O(N__753),
            .I(N__743));
    InMux I__73 (
            .O(N__750),
            .I(N__737));
    InMux I__72 (
            .O(N__749),
            .I(N__737));
    InMux I__71 (
            .O(N__746),
            .I(N__730));
    InMux I__70 (
            .O(N__743),
            .I(N__730));
    InMux I__69 (
            .O(N__742),
            .I(N__730));
    LocalMux I__68 (
            .O(N__737),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_3 ));
    LocalMux I__67 (
            .O(N__730),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_3 ));
    IoInMux I__66 (
            .O(N__725),
            .I(N__722));
    LocalMux I__65 (
            .O(N__722),
            .I(N__719));
    Span4Mux_s3_h I__64 (
            .O(N__719),
            .I(N__716));
    Odrv4 I__63 (
            .O(N__716),
            .I(RST_N_c_i));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_15_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB RST_N_ibuf_RNIBJGC_0 (
            .USERSIGNALTOGLOBALBUFFER(N__725),
            .GLOBALBUFFEROUTPUT(RST_N_c_i_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam RST_N_ibuf_RNIBJGC_LC_5_16_0.C_ON=1'b0;
    defparam RST_N_ibuf_RNIBJGC_LC_5_16_0.SEQ_MODE=4'b0000;
    defparam RST_N_ibuf_RNIBJGC_LC_5_16_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 RST_N_ibuf_RNIBJGC_LC_5_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1001),
            .lcout(RST_N_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counter_0_LC_11_13_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_0_LC_11_13_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter_0_LC_11_13_1 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \fsm_shiftRegs_inst1.counter_0_LC_11_13_1  (
            .in0(N__955),
            .in1(N__749),
            .in2(_gnd_net_),
            .in3(N__800),
            .lcout(\fsm_shiftRegs_inst1.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1423),
            .ce(),
            .sr(N__1385));
    defparam \fsm_shiftRegs_inst1.counter_1_LC_11_13_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_1_LC_11_13_2 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter_1_LC_11_13_2 .LUT_INIT=16'b1100010000001000;
    LogicCell40 \fsm_shiftRegs_inst1.counter_1_LC_11_13_2  (
            .in0(N__799),
            .in1(N__956),
            .in2(N__755),
            .in3(N__776),
            .lcout(\fsm_shiftRegs_inst1.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1423),
            .ce(),
            .sr(N__1385));
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_2_LC_12_13_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_2_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_2_LC_12_13_0 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \fsm_shiftRegs_inst1.counter_RNO_0_2_LC_12_13_0  (
            .in0(N__797),
            .in1(N__778),
            .in2(N__753),
            .in3(N__918),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counter_2_LC_12_13_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_2_LC_12_13_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter_2_LC_12_13_1 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \fsm_shiftRegs_inst1.counter_2_LC_12_13_1  (
            .in0(N__952),
            .in1(_gnd_net_),
            .in2(N__803),
            .in3(_gnd_net_),
            .lcout(\fsm_shiftRegs_inst1.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1426),
            .ce(),
            .sr(N__1388));
    defparam \fsm_shiftRegs_inst1.counter_RNIC589_1_LC_12_13_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_RNIC589_1_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.counter_RNIC589_1_LC_12_13_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \fsm_shiftRegs_inst1.counter_RNIC589_1_LC_12_13_3  (
            .in0(N__777),
            .in1(N__796),
            .in2(_gnd_net_),
            .in3(N__742),
            .lcout(\fsm_shiftRegs_inst1.N_123_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_3_LC_12_13_6 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_3_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_3_LC_12_13_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \fsm_shiftRegs_inst1.counter_RNO_0_3_LC_12_13_6  (
            .in0(N__798),
            .in1(N__779),
            .in2(N__754),
            .in3(N__919),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counter_3_LC_12_13_7 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_3_LC_12_13_7 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter_3_LC_12_13_7 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \fsm_shiftRegs_inst1.counter_3_LC_12_13_7  (
            .in0(N__953),
            .in1(_gnd_net_),
            .in2(N__758),
            .in3(_gnd_net_),
            .lcout(\fsm_shiftRegs_inst1.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1426),
            .ce(),
            .sr(N__1388));
    defparam \fsm_shiftRegs_inst1.current_state_1_LC_12_14_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_1_LC_12_14_2 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.current_state_1_LC_12_14_2 .LUT_INIT=16'b1111100011111010;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_1_LC_12_14_2  (
            .in0(N__954),
            .in1(N__920),
            .in2(N__1319),
            .in3(N__841),
            .lcout(\fsm_shiftRegs_inst1.current_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1424),
            .ce(),
            .sr(N__1386));
    defparam \fsm_shiftRegs_inst1.current_state_3_LC_12_14_7 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_3_LC_12_14_7 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.current_state_3_LC_12_14_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_3_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__1093),
            .in2(_gnd_net_),
            .in3(N__809),
            .lcout(\fsm_shiftRegs_inst1.current_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1424),
            .ce(),
            .sr(N__1386));
    defparam \fsm_shiftRegs_inst1.sel_stat_LC_12_15_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.sel_stat_LC_12_15_0 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.sel_stat_LC_12_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fsm_shiftRegs_inst1.sel_stat_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__893),
            .lcout(SELSTAT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1422),
            .ce(),
            .sr(N__1384));
    defparam \fsm_shiftRegs_inst1.sel_dyn_LC_12_15_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.sel_dyn_LC_12_15_2 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.sel_dyn_LC_12_15_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \fsm_shiftRegs_inst1.sel_dyn_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__1046),
            .in2(_gnd_net_),
            .in3(N__1208),
            .lcout(SELDYN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1422),
            .ce(),
            .sr(N__1384));
    defparam enableDin_aux_LC_13_11_2.C_ON=1'b0;
    defparam enableDin_aux_LC_13_11_2.SEQ_MODE=4'b1000;
    defparam enableDin_aux_LC_13_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 enableDin_aux_LC_13_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__854),
            .lcout(ENdin_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1433),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.en_fin_LC_13_12_6 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.en_fin_LC_13_12_6 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.en_fin_LC_13_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fsm_shiftRegs_inst1.en_fin_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1044),
            .lcout(enable_din),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1431),
            .ce(),
            .sr(N__1391));
    defparam \fsm_shiftRegs_inst1.counterDYN_RNO_0_3_LC_13_13_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counterDYN_RNO_0_3_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.counterDYN_RNO_0_3_LC_13_13_0 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \fsm_shiftRegs_inst1.counterDYN_RNO_0_3_LC_13_13_0  (
            .in0(N__825),
            .in1(N__1089),
            .in2(N__1067),
            .in3(N__1108),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counterDYN_3_LC_13_13_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counterDYN_3_LC_13_13_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counterDYN_3_LC_13_13_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fsm_shiftRegs_inst1.counterDYN_3_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__848),
            .in3(N__1039),
            .lcout(\fsm_shiftRegs_inst1.counterDYNZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1429),
            .ce(),
            .sr(N__1390));
    defparam \fsm_shiftRegs_inst1.counterDYN_0_LC_13_13_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counterDYN_0_LC_13_13_2 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counterDYN_0_LC_13_13_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \fsm_shiftRegs_inst1.counterDYN_0_LC_13_13_2  (
            .in0(N__1033),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1091),
            .lcout(\fsm_shiftRegs_inst1.counterDYNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1429),
            .ce(),
            .sr(N__1390));
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_2_LC_13_13_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_2_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_2_LC_13_13_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNO_0_2_LC_13_13_3  (
            .in0(N__1107),
            .in1(N__1064),
            .in2(N__1094),
            .in3(N__826),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_2_LC_13_13_4 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_2_LC_13_13_4 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.current_state_2_LC_13_13_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_2_LC_13_13_4  (
            .in0(N__1034),
            .in1(N__845),
            .in2(N__830),
            .in3(N__899),
            .lcout(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1429),
            .ce(),
            .sr(N__1390));
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_3_LC_13_13_5 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_3_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_3_LC_13_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNO_0_3_LC_13_13_5  (
            .in0(N__1106),
            .in1(N__1060),
            .in2(N__827),
            .in3(N__1032),
            .lcout(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counterDYN_2_LC_13_13_6 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counterDYN_2_LC_13_13_6 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counterDYN_2_LC_13_13_6 .LUT_INIT=16'b0111000010000000;
    LogicCell40 \fsm_shiftRegs_inst1.counterDYN_2_LC_13_13_6  (
            .in0(N__1065),
            .in1(N__1092),
            .in2(N__1045),
            .in3(N__1109),
            .lcout(\fsm_shiftRegs_inst1.counterDYNZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1429),
            .ce(),
            .sr(N__1390));
    defparam \fsm_shiftRegs_inst1.counterDYN_1_LC_13_13_7 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counterDYN_1_LC_13_13_7 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counterDYN_1_LC_13_13_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \fsm_shiftRegs_inst1.counterDYN_1_LC_13_13_7  (
            .in0(N__1090),
            .in1(N__1035),
            .in2(_gnd_net_),
            .in3(N__1066),
            .lcout(\fsm_shiftRegs_inst1.counterDYNZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1429),
            .ce(),
            .sr(N__1390));
    defparam \fsm_shiftRegs_inst1.signal_out_LC_13_14_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.signal_out_LC_13_14_0 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.signal_out_LC_13_14_0 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \fsm_shiftRegs_inst1.signal_out_LC_13_14_0  (
            .in0(N__1187),
            .in1(N__1361),
            .in2(N__1000),
            .in3(N__1043),
            .lcout(signal_out_fsm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1427),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_RNI7RPG_1_LC_13_14_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNI7RPG_1_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNI7RPG_1_LC_13_14_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNI7RPG_1_LC_13_14_2  (
            .in0(N__993),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__945),
            .lcout(\fsm_shiftRegs_inst1.un1_current_state4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_RNO_1_2_LC_13_14_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_1_2_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_1_2_LC_13_14_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNO_1_2_LC_13_14_3  (
            .in0(N__946),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__917),
            .lcout(\fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_4_LC_13_15_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_4_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_4_LC_13_15_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNO_0_4_LC_13_15_0  (
            .in0(N__1592),
            .in1(N__1234),
            .in2(N__1568),
            .in3(N__1531),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_4_LC_13_15_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_4_LC_13_15_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.current_state_4_LC_13_15_1 .LUT_INIT=16'b1100111011101110;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_4_LC_13_15_1  (
            .in0(N__1207),
            .in1(N__892),
            .in2(N__881),
            .in3(N__1217),
            .lcout(\fsm_shiftRegs_inst1.current_stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1425),
            .ce(),
            .sr(N__1387));
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_0_LC_13_15_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_0_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_0_LC_13_15_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNO_0_0_LC_13_15_2  (
            .in0(N__1564),
            .in1(N__1588),
            .in2(_gnd_net_),
            .in3(N__1530),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_0_LC_13_15_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_0_LC_13_15_3 .SEQ_MODE=4'b1011;
    defparam \fsm_shiftRegs_inst1.current_state_0_LC_13_15_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_0_LC_13_15_3  (
            .in0(N__1235),
            .in1(N__1206),
            .in2(N__878),
            .in3(N__1216),
            .lcout(\fsm_shiftRegs_inst1.current_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1425),
            .ce(),
            .sr(N__1387));
    defparam \fsm_shiftRegs_inst1.counter2_RNITAO81_7_LC_13_15_4 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter2_RNITAO81_7_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.counter2_RNITAO81_7_LC_13_15_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_RNITAO81_7_LC_13_15_4  (
            .in0(N__1510),
            .in1(N__1546),
            .in2(N__1496),
            .in3(N__1444),
            .lcout(\fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_RNIVA94_4_LC_13_15_5 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNIVA94_4_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNIVA94_4_LC_13_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNIVA94_4_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1205),
            .lcout(\fsm_shiftRegs_inst1.current_state_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.signal_aux_LC_13_15_7 .C_ON=1'b0;
    defparam \generator_inst1.signal_aux_LC_13_15_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.signal_aux_LC_13_15_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \generator_inst1.signal_aux_LC_13_15_7  (
            .in0(N__1186),
            .in1(N__1175),
            .in2(_gnd_net_),
            .in3(N__1169),
            .lcout(generated_signal_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1425),
            .ce(),
            .sr(N__1387));
    defparam \fsm_shiftRegs_inst1.bit_sequence_3_LC_14_13_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_3_LC_14_13_0 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_3_LC_14_13_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_3_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__1313),
            .in2(_gnd_net_),
            .in3(N__1139),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1432),
            .ce(N__1247),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_2_LC_14_13_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_2_LC_14_13_1 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_2_LC_14_13_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_2_LC_14_13_1  (
            .in0(N__1318),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1432),
            .ce(N__1247),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_4_LC_14_13_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_4_LC_14_13_2 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_4_LC_14_13_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_4_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(N__1314),
            .in2(_gnd_net_),
            .in3(N__1133),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1432),
            .ce(N__1247),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_6_LC_14_13_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_6_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_6_LC_14_13_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_6_LC_14_13_3  (
            .in0(N__1316),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1115),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1432),
            .ce(N__1247),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_7_LC_14_13_4 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_7_LC_14_13_4 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_7_LC_14_13_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_7_LC_14_13_4  (
            .in0(_gnd_net_),
            .in1(N__1317),
            .in2(_gnd_net_),
            .in3(N__1127),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1432),
            .ce(N__1247),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_5_LC_14_13_5 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_5_LC_14_13_5 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_5_LC_14_13_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_5_LC_14_13_5  (
            .in0(N__1315),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1121),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1432),
            .ce(N__1247),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_15_LC_14_14_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_15_LC_14_14_0 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_15_LC_14_14_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_15_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__1294),
            .in2(_gnd_net_),
            .in3(N__1331),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1430),
            .ce(N__1246),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_11_LC_14_14_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_11_LC_14_14_1 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_11_LC_14_14_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_11_LC_14_14_1  (
            .in0(N__1290),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1343),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1430),
            .ce(N__1246),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_12_LC_14_14_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_12_LC_14_14_2 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_12_LC_14_14_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_12_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__1291),
            .in2(_gnd_net_),
            .in3(N__1355),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1430),
            .ce(N__1246),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_13_LC_14_14_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_13_LC_14_14_3 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_13_LC_14_14_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_13_LC_14_14_3  (
            .in0(N__1292),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1349),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1430),
            .ce(N__1246),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_10_LC_14_14_4 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_10_LC_14_14_4 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_10_LC_14_14_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_10_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__1289),
            .in2(_gnd_net_),
            .in3(N__1325),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1430),
            .ce(N__1246),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_14_LC_14_14_5 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_14_LC_14_14_5 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_14_LC_14_14_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_14_LC_14_14_5  (
            .in0(N__1293),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1337),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1430),
            .ce(N__1246),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_9_LC_14_14_6 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_9_LC_14_14_6 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_9_LC_14_14_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_9_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__1296),
            .in2(_gnd_net_),
            .in3(N__1253),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1430),
            .ce(N__1246),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_8_LC_14_14_7 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_8_LC_14_14_7 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_8_LC_14_14_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_8_LC_14_14_7  (
            .in0(N__1295),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1259),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1430),
            .ce(N__1246),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counter2_0_LC_14_15_0 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_0_LC_14_15_0 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_0_LC_14_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_0_LC_14_15_0  (
            .in0(N__1475),
            .in1(N__1233),
            .in2(_gnd_net_),
            .in3(N__1220),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_0 ),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_0 ),
            .clk(N__1428),
            .ce(),
            .sr(N__1389));
    defparam \fsm_shiftRegs_inst1.counter2_1_LC_14_15_1 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_1_LC_14_15_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_1_LC_14_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_1_LC_14_15_1  (
            .in0(N__1471),
            .in1(N__1587),
            .in2(_gnd_net_),
            .in3(N__1571),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_1 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_0 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_1 ),
            .clk(N__1428),
            .ce(),
            .sr(N__1389));
    defparam \fsm_shiftRegs_inst1.counter2_2_LC_14_15_2 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_2_LC_14_15_2 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_2_LC_14_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_2_LC_14_15_2  (
            .in0(N__1476),
            .in1(N__1563),
            .in2(_gnd_net_),
            .in3(N__1550),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_2 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_1 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_2 ),
            .clk(N__1428),
            .ce(),
            .sr(N__1389));
    defparam \fsm_shiftRegs_inst1.counter2_3_LC_14_15_3 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_3_LC_14_15_3 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_3_LC_14_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_3_LC_14_15_3  (
            .in0(N__1472),
            .in1(N__1547),
            .in2(_gnd_net_),
            .in3(N__1535),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_3 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_2 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_3 ),
            .clk(N__1428),
            .ce(),
            .sr(N__1389));
    defparam \fsm_shiftRegs_inst1.counter2_4_LC_14_15_4 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_4_LC_14_15_4 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_4_LC_14_15_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_4_LC_14_15_4  (
            .in0(N__1477),
            .in1(_gnd_net_),
            .in2(N__1532),
            .in3(N__1514),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_4 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_3 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_4 ),
            .clk(N__1428),
            .ce(),
            .sr(N__1389));
    defparam \fsm_shiftRegs_inst1.counter2_5_LC_14_15_5 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_5_LC_14_15_5 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_5_LC_14_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_5_LC_14_15_5  (
            .in0(N__1473),
            .in1(N__1511),
            .in2(_gnd_net_),
            .in3(N__1499),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_5 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_4 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_5 ),
            .clk(N__1428),
            .ce(),
            .sr(N__1389));
    defparam \fsm_shiftRegs_inst1.counter2_6_LC_14_15_6 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_6_LC_14_15_6 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_6_LC_14_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_6_LC_14_15_6  (
            .in0(N__1478),
            .in1(N__1495),
            .in2(_gnd_net_),
            .in3(N__1481),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_6 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_5 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_6 ),
            .clk(N__1428),
            .ce(),
            .sr(N__1389));
    defparam \fsm_shiftRegs_inst1.counter2_7_LC_14_15_7 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter2_7_LC_14_15_7 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_7_LC_14_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_7_LC_14_15_7  (
            .in0(N__1474),
            .in1(N__1445),
            .in2(_gnd_net_),
            .in3(N__1448),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1428),
            .ce(),
            .sr(N__1389));
endmodule // top
