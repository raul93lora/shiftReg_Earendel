-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 20 2025 12:46:15

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    SDO_signal_out : out std_logic;
    RST_N : in std_logic;
    CLK_fast : in std_logic;
    CLK : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__6110\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \RST_N_c\ : std_logic;
signal \RST_N_c_i\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_21\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_72\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_28\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_70\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_71\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_20\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_26\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_27\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_69\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_25\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_24\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_22\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_23\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_66\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_67\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_68\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_64\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_65\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_83\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_13\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_29\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_30\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_12\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_11\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_10\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_63\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_14\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_12\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_13\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_73\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_84\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_82\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_74\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_75\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_14\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_31\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_32\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_33\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_1\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_81\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_19\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_7\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_62\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_2\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_8\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_9\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_61\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_10\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_11\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_8\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_9\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_6\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_7\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_5\ : std_logic;
signal \fsm_ctrl_inst1.un1_counter_statlt5_0_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_4\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_2\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_3\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_1\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_3\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_4\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_5\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_6\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_2\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_7\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_8\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_76\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_58\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_53\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_77\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_56\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_57\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_54\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_55\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_48\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_47\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_59\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_60\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_85\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_34\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_80\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_3\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_4\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_15\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_16\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_5\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_6\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_45\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_46\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_43\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_44\ : std_logic;
signal \bfn_6_21_0_\ : std_logic;
signal \fsm_ctrl_inst1.counter_stat_cry_0\ : std_logic;
signal \fsm_ctrl_inst1.counter_stat_cry_1\ : std_logic;
signal \fsm_ctrl_inst1.counter_stat_cry_2\ : std_logic;
signal \fsm_ctrl_inst1.counter_stat_cry_3\ : std_logic;
signal \fsm_ctrl_inst1.counter_stat_cry_4\ : std_logic;
signal \fsm_ctrl_inst1.current_state_i_1\ : std_logic;
signal \fsm_ctrl_inst1.counter_stat_cry_5\ : std_logic;
signal \fsm_ctrl_inst1.counter_state_0_i\ : std_logic;
signal \fsm_ctrl_inst1.counter_statZ0Z_3\ : std_logic;
signal \fsm_ctrl_inst1.counter_statZ0Z_1\ : std_logic;
signal \fsm_ctrl_inst1.counter_statZ0Z_6\ : std_logic;
signal \fsm_ctrl_inst1.counter_statZ0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.counter_statZ0Z_5\ : std_logic;
signal \fsm_ctrl_inst1.counter_statZ0Z_2\ : std_logic;
signal \fsm_ctrl_inst1.current_state_ns_i_a3_0_4_1_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.counter_statZ0Z_4\ : std_logic;
signal \fsm_ctrl_inst1.current_state_ns_i_a3_0_5_1_cascade_\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_0\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_1\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_9\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_10\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_11\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_12\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_13\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_14\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSR_cnvZ0Z_0\ : std_logic;
signal \toggle_clk_uC4_0\ : std_logic;
signal \fsm_ctrl_inst1_CLK_uC_1_i\ : std_logic;
signal \STATSR_cnv_0\ : std_logic;
signal \fsm_ctrl_inst1.counter_idlelde_0_a3_0_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_78\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_79\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_52\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_35\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_49\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_36\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_37\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_50\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_51\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_38\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_39\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_86\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_17\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_18\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_42\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_40\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_41\ : std_logic;
signal \fsm_ctrl_inst1.current_state_i_g_0\ : std_logic;
signal \fsm_ctrl_inst1.current_state_i_0\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_15\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_87\ : std_logic;
signal \fsm_ctrl_inst1.N_119_0\ : std_logic;
signal \fsm_ctrl_inst1.N_105_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.counter_dinZ0Z_3\ : std_logic;
signal \fsm_ctrl_inst1.counter_dinZ0Z_2\ : std_logic;
signal \fsm_ctrl_inst1.counter_dinZ0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.counter_dinZ0Z_1\ : std_logic;
signal \SEL_REG\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_15\ : std_logic;
signal \SDO_signal_out_c\ : std_logic;
signal \fsm_ctrl_inst1.current_state_ns_0_i_0_1_0\ : std_logic;
signal \fsm_ctrl_inst1.N_122_2\ : std_logic;
signal \fsm_ctrl_inst1.counter_idleZ0Z_0\ : std_logic;
signal \bfn_7_25_0_\ : std_logic;
signal \fsm_ctrl_inst1.counter_idleZ0Z_1\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_cry_0\ : std_logic;
signal \fsm_ctrl_inst1.counter_idleZ0Z_2\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_cry_1\ : std_logic;
signal \fsm_ctrl_inst1.counter_idleZ0Z_3\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_cry_2\ : std_logic;
signal \fsm_ctrl_inst1.current_state_23_d_i\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_cry_3\ : std_logic;
signal \fsm_ctrl_inst1.counter_idleZ0Z_4\ : std_logic;
signal \fsm_ctrl_inst1.counter_idlee_0_i\ : std_logic;
signal \fsm_ctrl_inst1.toggle_clk_uC3Z0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.toggle_clk_uC2Z0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.current_stateZ0Z_1\ : std_logic;
signal \fsm_ctrl_inst1.current_stateZ0Z_0\ : std_logic;
signal \CLK_c_g\ : std_logic;
signal \fsm_ctrl_inst1.toggle_clk_uCZ0Z1\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_87\ : std_logic;
signal \MOSI\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_85\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_86\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_0\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_3\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_1\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_2\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_84\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_83\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_4\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_5\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_82\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_6\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_7\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_8\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_9\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_10\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_11\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_79\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_80\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_81\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_78\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_77\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_14\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_12\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_13\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_15\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_74\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_75\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_76\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_73\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_16\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_71\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_72\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_68\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_69\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_70\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_66\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_67\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_65\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_62\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_61\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_63\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_64\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_17\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_18\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_56\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_60\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_57\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_58\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_59\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_50\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_49\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_53\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_54\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_55\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_51\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_52\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_19\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_20\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_33\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_34\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_21\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_30\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_22\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_23\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_31\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_32\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_24\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_25\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_26\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_29\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_27\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_28\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_48\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_42\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_43\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_44\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_45\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_46\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_47\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_41\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_40\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_38\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_39\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_35\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_36\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_37\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \CLK_fast_0_c_g\ : std_logic;
signal \N_224_g\ : std_logic;
signal \RST_N_c_i_g\ : std_logic;

signal \CLK_fast_wire\ : std_logic;
signal \CLK_wire\ : std_logic;
signal \RST_N_wire\ : std_logic;
signal \SDO_signal_out_wire\ : std_logic;

begin
    \CLK_fast_wire\ <= CLK_fast;
    \CLK_wire\ <= CLK;
    \RST_N_wire\ <= RST_N;
    SDO_signal_out <= \SDO_signal_out_wire\;

    \CLK_fast_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6108\,
            GLOBALBUFFEROUTPUT => \CLK_fast_0_c_g\
        );

    \CLK_fast_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6110\,
            DIN => \N__6109\,
            DOUT => \N__6108\,
            PACKAGEPIN => \CLK_fast_wire\
        );

    \CLK_fast_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6110\,
            PADOUT => \N__6109\,
            PADIN => \N__6108\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6098\,
            GLOBALBUFFEROUTPUT => \CLK_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6100\,
            DIN => \N__6099\,
            DOUT => \N__6098\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6100\,
            PADOUT => \N__6099\,
            PADIN => \N__6098\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RST_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6089\,
            DIN => \N__6088\,
            DOUT => \N__6087\,
            PACKAGEPIN => \RST_N_wire\
        );

    \RST_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6089\,
            PADOUT => \N__6088\,
            PADIN => \N__6087\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RST_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SDO_signal_out_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6080\,
            DIN => \N__6079\,
            DOUT => \N__6078\,
            PACKAGEPIN => \SDO_signal_out_wire\
        );

    \SDO_signal_out_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6080\,
            PADOUT => \N__6079\,
            PADIN => \N__6078\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4204\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1255\ : InMux
    port map (
            O => \N__6061\,
            I => \N__6058\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6058\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_44\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6055\,
            I => \N__6052\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__6052\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_45\
        );

    \I__1251\ : InMux
    port map (
            O => \N__6049\,
            I => \N__6046\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__6046\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_46\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6043\,
            I => \N__6040\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6040\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_47\
        );

    \I__1247\ : InMux
    port map (
            O => \N__6037\,
            I => \N__6034\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__6034\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_41\
        );

    \I__1245\ : InMux
    port map (
            O => \N__6031\,
            I => \N__6028\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__6028\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_40\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6025\,
            I => \N__6022\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__6022\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_38\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6019\,
            I => \N__6016\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__6016\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_39\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6013\,
            I => \N__6010\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6010\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_35\
        );

    \I__1237\ : InMux
    port map (
            O => \N__6007\,
            I => \N__6004\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__6004\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_36\
        );

    \I__1235\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5998\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__5998\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_37\
        );

    \I__1233\ : ClkMux
    port map (
            O => \N__5995\,
            I => \N__5902\
        );

    \I__1232\ : ClkMux
    port map (
            O => \N__5994\,
            I => \N__5902\
        );

    \I__1231\ : ClkMux
    port map (
            O => \N__5993\,
            I => \N__5902\
        );

    \I__1230\ : ClkMux
    port map (
            O => \N__5992\,
            I => \N__5902\
        );

    \I__1229\ : ClkMux
    port map (
            O => \N__5991\,
            I => \N__5902\
        );

    \I__1228\ : ClkMux
    port map (
            O => \N__5990\,
            I => \N__5902\
        );

    \I__1227\ : ClkMux
    port map (
            O => \N__5989\,
            I => \N__5902\
        );

    \I__1226\ : ClkMux
    port map (
            O => \N__5988\,
            I => \N__5902\
        );

    \I__1225\ : ClkMux
    port map (
            O => \N__5987\,
            I => \N__5902\
        );

    \I__1224\ : ClkMux
    port map (
            O => \N__5986\,
            I => \N__5902\
        );

    \I__1223\ : ClkMux
    port map (
            O => \N__5985\,
            I => \N__5902\
        );

    \I__1222\ : ClkMux
    port map (
            O => \N__5984\,
            I => \N__5902\
        );

    \I__1221\ : ClkMux
    port map (
            O => \N__5983\,
            I => \N__5902\
        );

    \I__1220\ : ClkMux
    port map (
            O => \N__5982\,
            I => \N__5902\
        );

    \I__1219\ : ClkMux
    port map (
            O => \N__5981\,
            I => \N__5902\
        );

    \I__1218\ : ClkMux
    port map (
            O => \N__5980\,
            I => \N__5902\
        );

    \I__1217\ : ClkMux
    port map (
            O => \N__5979\,
            I => \N__5902\
        );

    \I__1216\ : ClkMux
    port map (
            O => \N__5978\,
            I => \N__5902\
        );

    \I__1215\ : ClkMux
    port map (
            O => \N__5977\,
            I => \N__5902\
        );

    \I__1214\ : ClkMux
    port map (
            O => \N__5976\,
            I => \N__5902\
        );

    \I__1213\ : ClkMux
    port map (
            O => \N__5975\,
            I => \N__5902\
        );

    \I__1212\ : ClkMux
    port map (
            O => \N__5974\,
            I => \N__5902\
        );

    \I__1211\ : ClkMux
    port map (
            O => \N__5973\,
            I => \N__5902\
        );

    \I__1210\ : ClkMux
    port map (
            O => \N__5972\,
            I => \N__5902\
        );

    \I__1209\ : ClkMux
    port map (
            O => \N__5971\,
            I => \N__5902\
        );

    \I__1208\ : ClkMux
    port map (
            O => \N__5970\,
            I => \N__5902\
        );

    \I__1207\ : ClkMux
    port map (
            O => \N__5969\,
            I => \N__5902\
        );

    \I__1206\ : ClkMux
    port map (
            O => \N__5968\,
            I => \N__5902\
        );

    \I__1205\ : ClkMux
    port map (
            O => \N__5967\,
            I => \N__5902\
        );

    \I__1204\ : ClkMux
    port map (
            O => \N__5966\,
            I => \N__5902\
        );

    \I__1203\ : ClkMux
    port map (
            O => \N__5965\,
            I => \N__5902\
        );

    \I__1202\ : GlobalMux
    port map (
            O => \N__5902\,
            I => \N__5899\
        );

    \I__1201\ : gio2CtrlBuf
    port map (
            O => \N__5899\,
            I => \CLK_fast_0_c_g\
        );

    \I__1200\ : CEMux
    port map (
            O => \N__5896\,
            I => \N__5818\
        );

    \I__1199\ : CEMux
    port map (
            O => \N__5895\,
            I => \N__5818\
        );

    \I__1198\ : CEMux
    port map (
            O => \N__5894\,
            I => \N__5818\
        );

    \I__1197\ : CEMux
    port map (
            O => \N__5893\,
            I => \N__5818\
        );

    \I__1196\ : CEMux
    port map (
            O => \N__5892\,
            I => \N__5818\
        );

    \I__1195\ : CEMux
    port map (
            O => \N__5891\,
            I => \N__5818\
        );

    \I__1194\ : CEMux
    port map (
            O => \N__5890\,
            I => \N__5818\
        );

    \I__1193\ : CEMux
    port map (
            O => \N__5889\,
            I => \N__5818\
        );

    \I__1192\ : CEMux
    port map (
            O => \N__5888\,
            I => \N__5818\
        );

    \I__1191\ : CEMux
    port map (
            O => \N__5887\,
            I => \N__5818\
        );

    \I__1190\ : CEMux
    port map (
            O => \N__5886\,
            I => \N__5818\
        );

    \I__1189\ : CEMux
    port map (
            O => \N__5885\,
            I => \N__5818\
        );

    \I__1188\ : CEMux
    port map (
            O => \N__5884\,
            I => \N__5818\
        );

    \I__1187\ : CEMux
    port map (
            O => \N__5883\,
            I => \N__5818\
        );

    \I__1186\ : CEMux
    port map (
            O => \N__5882\,
            I => \N__5818\
        );

    \I__1185\ : CEMux
    port map (
            O => \N__5881\,
            I => \N__5818\
        );

    \I__1184\ : CEMux
    port map (
            O => \N__5880\,
            I => \N__5818\
        );

    \I__1183\ : CEMux
    port map (
            O => \N__5879\,
            I => \N__5818\
        );

    \I__1182\ : CEMux
    port map (
            O => \N__5878\,
            I => \N__5818\
        );

    \I__1181\ : CEMux
    port map (
            O => \N__5877\,
            I => \N__5818\
        );

    \I__1180\ : CEMux
    port map (
            O => \N__5876\,
            I => \N__5818\
        );

    \I__1179\ : CEMux
    port map (
            O => \N__5875\,
            I => \N__5818\
        );

    \I__1178\ : CEMux
    port map (
            O => \N__5874\,
            I => \N__5818\
        );

    \I__1177\ : CEMux
    port map (
            O => \N__5873\,
            I => \N__5818\
        );

    \I__1176\ : CEMux
    port map (
            O => \N__5872\,
            I => \N__5818\
        );

    \I__1175\ : CEMux
    port map (
            O => \N__5871\,
            I => \N__5818\
        );

    \I__1174\ : GlobalMux
    port map (
            O => \N__5818\,
            I => \N__5815\
        );

    \I__1173\ : gio2CtrlBuf
    port map (
            O => \N__5815\,
            I => \N_224_g\
        );

    \I__1172\ : SRMux
    port map (
            O => \N__5812\,
            I => \N__5635\
        );

    \I__1171\ : SRMux
    port map (
            O => \N__5811\,
            I => \N__5635\
        );

    \I__1170\ : SRMux
    port map (
            O => \N__5810\,
            I => \N__5635\
        );

    \I__1169\ : SRMux
    port map (
            O => \N__5809\,
            I => \N__5635\
        );

    \I__1168\ : SRMux
    port map (
            O => \N__5808\,
            I => \N__5635\
        );

    \I__1167\ : SRMux
    port map (
            O => \N__5807\,
            I => \N__5635\
        );

    \I__1166\ : SRMux
    port map (
            O => \N__5806\,
            I => \N__5635\
        );

    \I__1165\ : SRMux
    port map (
            O => \N__5805\,
            I => \N__5635\
        );

    \I__1164\ : SRMux
    port map (
            O => \N__5804\,
            I => \N__5635\
        );

    \I__1163\ : SRMux
    port map (
            O => \N__5803\,
            I => \N__5635\
        );

    \I__1162\ : SRMux
    port map (
            O => \N__5802\,
            I => \N__5635\
        );

    \I__1161\ : SRMux
    port map (
            O => \N__5801\,
            I => \N__5635\
        );

    \I__1160\ : SRMux
    port map (
            O => \N__5800\,
            I => \N__5635\
        );

    \I__1159\ : SRMux
    port map (
            O => \N__5799\,
            I => \N__5635\
        );

    \I__1158\ : SRMux
    port map (
            O => \N__5798\,
            I => \N__5635\
        );

    \I__1157\ : SRMux
    port map (
            O => \N__5797\,
            I => \N__5635\
        );

    \I__1156\ : SRMux
    port map (
            O => \N__5796\,
            I => \N__5635\
        );

    \I__1155\ : SRMux
    port map (
            O => \N__5795\,
            I => \N__5635\
        );

    \I__1154\ : SRMux
    port map (
            O => \N__5794\,
            I => \N__5635\
        );

    \I__1153\ : SRMux
    port map (
            O => \N__5793\,
            I => \N__5635\
        );

    \I__1152\ : SRMux
    port map (
            O => \N__5792\,
            I => \N__5635\
        );

    \I__1151\ : SRMux
    port map (
            O => \N__5791\,
            I => \N__5635\
        );

    \I__1150\ : SRMux
    port map (
            O => \N__5790\,
            I => \N__5635\
        );

    \I__1149\ : SRMux
    port map (
            O => \N__5789\,
            I => \N__5635\
        );

    \I__1148\ : SRMux
    port map (
            O => \N__5788\,
            I => \N__5635\
        );

    \I__1147\ : SRMux
    port map (
            O => \N__5787\,
            I => \N__5635\
        );

    \I__1146\ : SRMux
    port map (
            O => \N__5786\,
            I => \N__5635\
        );

    \I__1145\ : SRMux
    port map (
            O => \N__5785\,
            I => \N__5635\
        );

    \I__1144\ : SRMux
    port map (
            O => \N__5784\,
            I => \N__5635\
        );

    \I__1143\ : SRMux
    port map (
            O => \N__5783\,
            I => \N__5635\
        );

    \I__1142\ : SRMux
    port map (
            O => \N__5782\,
            I => \N__5635\
        );

    \I__1141\ : SRMux
    port map (
            O => \N__5781\,
            I => \N__5635\
        );

    \I__1140\ : SRMux
    port map (
            O => \N__5780\,
            I => \N__5635\
        );

    \I__1139\ : SRMux
    port map (
            O => \N__5779\,
            I => \N__5635\
        );

    \I__1138\ : SRMux
    port map (
            O => \N__5778\,
            I => \N__5635\
        );

    \I__1137\ : SRMux
    port map (
            O => \N__5777\,
            I => \N__5635\
        );

    \I__1136\ : SRMux
    port map (
            O => \N__5776\,
            I => \N__5635\
        );

    \I__1135\ : SRMux
    port map (
            O => \N__5775\,
            I => \N__5635\
        );

    \I__1134\ : SRMux
    port map (
            O => \N__5774\,
            I => \N__5635\
        );

    \I__1133\ : SRMux
    port map (
            O => \N__5773\,
            I => \N__5635\
        );

    \I__1132\ : SRMux
    port map (
            O => \N__5772\,
            I => \N__5635\
        );

    \I__1131\ : SRMux
    port map (
            O => \N__5771\,
            I => \N__5635\
        );

    \I__1130\ : SRMux
    port map (
            O => \N__5770\,
            I => \N__5635\
        );

    \I__1129\ : SRMux
    port map (
            O => \N__5769\,
            I => \N__5635\
        );

    \I__1128\ : SRMux
    port map (
            O => \N__5768\,
            I => \N__5635\
        );

    \I__1127\ : SRMux
    port map (
            O => \N__5767\,
            I => \N__5635\
        );

    \I__1126\ : SRMux
    port map (
            O => \N__5766\,
            I => \N__5635\
        );

    \I__1125\ : SRMux
    port map (
            O => \N__5765\,
            I => \N__5635\
        );

    \I__1124\ : SRMux
    port map (
            O => \N__5764\,
            I => \N__5635\
        );

    \I__1123\ : SRMux
    port map (
            O => \N__5763\,
            I => \N__5635\
        );

    \I__1122\ : SRMux
    port map (
            O => \N__5762\,
            I => \N__5635\
        );

    \I__1121\ : SRMux
    port map (
            O => \N__5761\,
            I => \N__5635\
        );

    \I__1120\ : SRMux
    port map (
            O => \N__5760\,
            I => \N__5635\
        );

    \I__1119\ : SRMux
    port map (
            O => \N__5759\,
            I => \N__5635\
        );

    \I__1118\ : SRMux
    port map (
            O => \N__5758\,
            I => \N__5635\
        );

    \I__1117\ : SRMux
    port map (
            O => \N__5757\,
            I => \N__5635\
        );

    \I__1116\ : SRMux
    port map (
            O => \N__5756\,
            I => \N__5635\
        );

    \I__1115\ : SRMux
    port map (
            O => \N__5755\,
            I => \N__5635\
        );

    \I__1114\ : SRMux
    port map (
            O => \N__5754\,
            I => \N__5635\
        );

    \I__1113\ : GlobalMux
    port map (
            O => \N__5635\,
            I => \N__5632\
        );

    \I__1112\ : gio2CtrlBuf
    port map (
            O => \N__5632\,
            I => \RST_N_c_i_g\
        );

    \I__1111\ : InMux
    port map (
            O => \N__5629\,
            I => \N__5626\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__5626\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_25\
        );

    \I__1109\ : InMux
    port map (
            O => \N__5623\,
            I => \N__5620\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__5620\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_26\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5614\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__5614\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_29\
        );

    \I__1105\ : InMux
    port map (
            O => \N__5611\,
            I => \N__5608\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5608\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_27\
        );

    \I__1103\ : InMux
    port map (
            O => \N__5605\,
            I => \N__5602\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5602\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_28\
        );

    \I__1101\ : InMux
    port map (
            O => \N__5599\,
            I => \N__5596\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__5596\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_48\
        );

    \I__1099\ : InMux
    port map (
            O => \N__5593\,
            I => \N__5590\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__5590\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_42\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5587\,
            I => \N__5584\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__5584\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_43\
        );

    \I__1095\ : InMux
    port map (
            O => \N__5581\,
            I => \N__5578\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__5578\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_33\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5575\,
            I => \N__5572\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__5572\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_34\
        );

    \I__1091\ : InMux
    port map (
            O => \N__5569\,
            I => \N__5566\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__5566\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_21\
        );

    \I__1089\ : InMux
    port map (
            O => \N__5563\,
            I => \N__5560\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__5560\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_30\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5554\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5554\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_22\
        );

    \I__1085\ : InMux
    port map (
            O => \N__5551\,
            I => \N__5548\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__5548\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_23\
        );

    \I__1083\ : InMux
    port map (
            O => \N__5545\,
            I => \N__5542\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__5542\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_31\
        );

    \I__1081\ : InMux
    port map (
            O => \N__5539\,
            I => \N__5536\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__5536\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_32\
        );

    \I__1079\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5530\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__5530\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_24\
        );

    \I__1077\ : InMux
    port map (
            O => \N__5527\,
            I => \N__5524\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5524\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_50\
        );

    \I__1075\ : InMux
    port map (
            O => \N__5521\,
            I => \N__5518\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__5518\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_49\
        );

    \I__1073\ : InMux
    port map (
            O => \N__5515\,
            I => \N__5512\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__5512\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_53\
        );

    \I__1071\ : InMux
    port map (
            O => \N__5509\,
            I => \N__5506\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__5506\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_54\
        );

    \I__1069\ : InMux
    port map (
            O => \N__5503\,
            I => \N__5500\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__5500\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_55\
        );

    \I__1067\ : InMux
    port map (
            O => \N__5497\,
            I => \N__5494\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__5494\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_51\
        );

    \I__1065\ : InMux
    port map (
            O => \N__5491\,
            I => \N__5488\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__5488\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_52\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5485\,
            I => \N__5482\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__5482\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_19\
        );

    \I__1061\ : InMux
    port map (
            O => \N__5479\,
            I => \N__5476\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__5476\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_20\
        );

    \I__1059\ : InMux
    port map (
            O => \N__5473\,
            I => \N__5470\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__5470\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_61\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5467\,
            I => \N__5464\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__5464\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_63\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5461\,
            I => \N__5458\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__5458\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_64\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5452\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__5452\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_17\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5449\,
            I => \N__5446\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__5446\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_18\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5440\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__5440\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_56\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5437\,
            I => \N__5434\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__5434\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_60\
        );

    \I__1045\ : InMux
    port map (
            O => \N__5431\,
            I => \N__5428\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__5428\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_57\
        );

    \I__1043\ : InMux
    port map (
            O => \N__5425\,
            I => \N__5422\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__5422\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_58\
        );

    \I__1041\ : InMux
    port map (
            O => \N__5419\,
            I => \N__5416\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__5416\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_59\
        );

    \I__1039\ : InMux
    port map (
            O => \N__5413\,
            I => \N__5410\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__5410\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_71\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5407\,
            I => \N__5404\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__5404\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_72\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5401\,
            I => \N__5398\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__5398\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_68\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5392\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__5392\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_69\
        );

    \I__1031\ : InMux
    port map (
            O => \N__5389\,
            I => \N__5386\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__5386\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_70\
        );

    \I__1029\ : InMux
    port map (
            O => \N__5383\,
            I => \N__5380\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__5380\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_66\
        );

    \I__1027\ : InMux
    port map (
            O => \N__5377\,
            I => \N__5374\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__5374\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_67\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5371\,
            I => \N__5368\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__5368\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_65\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5365\,
            I => \N__5362\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__5362\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_62\
        );

    \I__1021\ : InMux
    port map (
            O => \N__5359\,
            I => \N__5356\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__5356\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_14\
        );

    \I__1019\ : InMux
    port map (
            O => \N__5353\,
            I => \N__5350\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5350\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_12\
        );

    \I__1017\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5344\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__5344\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_13\
        );

    \I__1015\ : InMux
    port map (
            O => \N__5341\,
            I => \N__5338\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5338\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_15\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5335\,
            I => \N__5332\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5332\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_74\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5329\,
            I => \N__5326\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__5326\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_75\
        );

    \I__1009\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5320\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5320\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_76\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5317\,
            I => \N__5314\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__5314\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_73\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5311\,
            I => \N__5308\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__5308\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_16\
        );

    \I__1003\ : InMux
    port map (
            O => \N__5305\,
            I => \N__5302\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__5302\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_8\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5299\,
            I => \N__5296\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__5296\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_9\
        );

    \I__999\ : InMux
    port map (
            O => \N__5293\,
            I => \N__5290\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__5290\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_10\
        );

    \I__997\ : InMux
    port map (
            O => \N__5287\,
            I => \N__5284\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5284\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_11\
        );

    \I__995\ : InMux
    port map (
            O => \N__5281\,
            I => \N__5278\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5278\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_79\
        );

    \I__993\ : InMux
    port map (
            O => \N__5275\,
            I => \N__5272\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__5272\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_80\
        );

    \I__991\ : InMux
    port map (
            O => \N__5269\,
            I => \N__5266\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__5266\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_81\
        );

    \I__989\ : InMux
    port map (
            O => \N__5263\,
            I => \N__5260\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__5260\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_78\
        );

    \I__987\ : InMux
    port map (
            O => \N__5257\,
            I => \N__5254\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__5254\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_77\
        );

    \I__985\ : InMux
    port map (
            O => \N__5251\,
            I => \N__5248\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__5248\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_1\
        );

    \I__983\ : InMux
    port map (
            O => \N__5245\,
            I => \N__5242\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5242\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_2\
        );

    \I__981\ : InMux
    port map (
            O => \N__5239\,
            I => \N__5236\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__5236\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_84\
        );

    \I__979\ : InMux
    port map (
            O => \N__5233\,
            I => \N__5230\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5230\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_83\
        );

    \I__977\ : InMux
    port map (
            O => \N__5227\,
            I => \N__5224\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__5224\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_4\
        );

    \I__975\ : InMux
    port map (
            O => \N__5221\,
            I => \N__5218\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__5218\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_5\
        );

    \I__973\ : InMux
    port map (
            O => \N__5215\,
            I => \N__5212\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__5212\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_82\
        );

    \I__971\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5206\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__5206\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_6\
        );

    \I__969\ : InMux
    port map (
            O => \N__5203\,
            I => \N__5200\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5200\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_7\
        );

    \I__967\ : InMux
    port map (
            O => \N__5197\,
            I => \N__5194\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5194\,
            I => \fsm_ctrl_inst1.toggle_clk_uC2Z0Z_0\
        );

    \I__965\ : InMux
    port map (
            O => \N__5191\,
            I => \N__5162\
        );

    \I__964\ : InMux
    port map (
            O => \N__5190\,
            I => \N__5155\
        );

    \I__963\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5155\
        );

    \I__962\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5155\
        );

    \I__961\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5146\
        );

    \I__960\ : InMux
    port map (
            O => \N__5186\,
            I => \N__5146\
        );

    \I__959\ : InMux
    port map (
            O => \N__5185\,
            I => \N__5146\
        );

    \I__958\ : InMux
    port map (
            O => \N__5184\,
            I => \N__5146\
        );

    \I__957\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5139\
        );

    \I__956\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5139\
        );

    \I__955\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5139\
        );

    \I__954\ : InMux
    port map (
            O => \N__5180\,
            I => \N__5128\
        );

    \I__953\ : InMux
    port map (
            O => \N__5179\,
            I => \N__5128\
        );

    \I__952\ : InMux
    port map (
            O => \N__5178\,
            I => \N__5128\
        );

    \I__951\ : InMux
    port map (
            O => \N__5177\,
            I => \N__5128\
        );

    \I__950\ : InMux
    port map (
            O => \N__5176\,
            I => \N__5128\
        );

    \I__949\ : InMux
    port map (
            O => \N__5175\,
            I => \N__5119\
        );

    \I__948\ : InMux
    port map (
            O => \N__5174\,
            I => \N__5119\
        );

    \I__947\ : InMux
    port map (
            O => \N__5173\,
            I => \N__5119\
        );

    \I__946\ : InMux
    port map (
            O => \N__5172\,
            I => \N__5119\
        );

    \I__945\ : InMux
    port map (
            O => \N__5171\,
            I => \N__5095\
        );

    \I__944\ : InMux
    port map (
            O => \N__5170\,
            I => \N__5090\
        );

    \I__943\ : InMux
    port map (
            O => \N__5169\,
            I => \N__5090\
        );

    \I__942\ : InMux
    port map (
            O => \N__5168\,
            I => \N__5045\
        );

    \I__941\ : InMux
    port map (
            O => \N__5167\,
            I => \N__5040\
        );

    \I__940\ : InMux
    port map (
            O => \N__5166\,
            I => \N__5040\
        );

    \I__939\ : InMux
    port map (
            O => \N__5165\,
            I => \N__5037\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5162\,
            I => \N__5030\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__5155\,
            I => \N__5025\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__5146\,
            I => \N__5025\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__5139\,
            I => \N__5022\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5128\,
            I => \N__5017\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__5119\,
            I => \N__5017\
        );

    \I__932\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5012\
        );

    \I__931\ : InMux
    port map (
            O => \N__5117\,
            I => \N__5012\
        );

    \I__930\ : InMux
    port map (
            O => \N__5116\,
            I => \N__4999\
        );

    \I__929\ : InMux
    port map (
            O => \N__5115\,
            I => \N__4999\
        );

    \I__928\ : InMux
    port map (
            O => \N__5114\,
            I => \N__4999\
        );

    \I__927\ : InMux
    port map (
            O => \N__5113\,
            I => \N__4999\
        );

    \I__926\ : InMux
    port map (
            O => \N__5112\,
            I => \N__4999\
        );

    \I__925\ : InMux
    port map (
            O => \N__5111\,
            I => \N__4999\
        );

    \I__924\ : InMux
    port map (
            O => \N__5110\,
            I => \N__4986\
        );

    \I__923\ : InMux
    port map (
            O => \N__5109\,
            I => \N__4986\
        );

    \I__922\ : InMux
    port map (
            O => \N__5108\,
            I => \N__4986\
        );

    \I__921\ : InMux
    port map (
            O => \N__5107\,
            I => \N__4986\
        );

    \I__920\ : InMux
    port map (
            O => \N__5106\,
            I => \N__4986\
        );

    \I__919\ : InMux
    port map (
            O => \N__5105\,
            I => \N__4986\
        );

    \I__918\ : InMux
    port map (
            O => \N__5104\,
            I => \N__4971\
        );

    \I__917\ : InMux
    port map (
            O => \N__5103\,
            I => \N__4971\
        );

    \I__916\ : InMux
    port map (
            O => \N__5102\,
            I => \N__4971\
        );

    \I__915\ : InMux
    port map (
            O => \N__5101\,
            I => \N__4971\
        );

    \I__914\ : InMux
    port map (
            O => \N__5100\,
            I => \N__4971\
        );

    \I__913\ : InMux
    port map (
            O => \N__5099\,
            I => \N__4971\
        );

    \I__912\ : InMux
    port map (
            O => \N__5098\,
            I => \N__4971\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__5095\,
            I => \N__4966\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__5090\,
            I => \N__4966\
        );

    \I__909\ : InMux
    port map (
            O => \N__5089\,
            I => \N__4949\
        );

    \I__908\ : InMux
    port map (
            O => \N__5088\,
            I => \N__4949\
        );

    \I__907\ : InMux
    port map (
            O => \N__5087\,
            I => \N__4949\
        );

    \I__906\ : InMux
    port map (
            O => \N__5086\,
            I => \N__4949\
        );

    \I__905\ : InMux
    port map (
            O => \N__5085\,
            I => \N__4949\
        );

    \I__904\ : InMux
    port map (
            O => \N__5084\,
            I => \N__4949\
        );

    \I__903\ : InMux
    port map (
            O => \N__5083\,
            I => \N__4949\
        );

    \I__902\ : InMux
    port map (
            O => \N__5082\,
            I => \N__4949\
        );

    \I__901\ : InMux
    port map (
            O => \N__5081\,
            I => \N__4932\
        );

    \I__900\ : InMux
    port map (
            O => \N__5080\,
            I => \N__4932\
        );

    \I__899\ : InMux
    port map (
            O => \N__5079\,
            I => \N__4932\
        );

    \I__898\ : InMux
    port map (
            O => \N__5078\,
            I => \N__4932\
        );

    \I__897\ : InMux
    port map (
            O => \N__5077\,
            I => \N__4932\
        );

    \I__896\ : InMux
    port map (
            O => \N__5076\,
            I => \N__4932\
        );

    \I__895\ : InMux
    port map (
            O => \N__5075\,
            I => \N__4932\
        );

    \I__894\ : InMux
    port map (
            O => \N__5074\,
            I => \N__4932\
        );

    \I__893\ : InMux
    port map (
            O => \N__5073\,
            I => \N__4915\
        );

    \I__892\ : InMux
    port map (
            O => \N__5072\,
            I => \N__4915\
        );

    \I__891\ : InMux
    port map (
            O => \N__5071\,
            I => \N__4915\
        );

    \I__890\ : InMux
    port map (
            O => \N__5070\,
            I => \N__4915\
        );

    \I__889\ : InMux
    port map (
            O => \N__5069\,
            I => \N__4915\
        );

    \I__888\ : InMux
    port map (
            O => \N__5068\,
            I => \N__4915\
        );

    \I__887\ : InMux
    port map (
            O => \N__5067\,
            I => \N__4915\
        );

    \I__886\ : InMux
    port map (
            O => \N__5066\,
            I => \N__4915\
        );

    \I__885\ : InMux
    port map (
            O => \N__5065\,
            I => \N__4898\
        );

    \I__884\ : InMux
    port map (
            O => \N__5064\,
            I => \N__4898\
        );

    \I__883\ : InMux
    port map (
            O => \N__5063\,
            I => \N__4898\
        );

    \I__882\ : InMux
    port map (
            O => \N__5062\,
            I => \N__4898\
        );

    \I__881\ : InMux
    port map (
            O => \N__5061\,
            I => \N__4898\
        );

    \I__880\ : InMux
    port map (
            O => \N__5060\,
            I => \N__4898\
        );

    \I__879\ : InMux
    port map (
            O => \N__5059\,
            I => \N__4898\
        );

    \I__878\ : InMux
    port map (
            O => \N__5058\,
            I => \N__4898\
        );

    \I__877\ : InMux
    port map (
            O => \N__5057\,
            I => \N__4895\
        );

    \I__876\ : InMux
    port map (
            O => \N__5056\,
            I => \N__4878\
        );

    \I__875\ : InMux
    port map (
            O => \N__5055\,
            I => \N__4878\
        );

    \I__874\ : InMux
    port map (
            O => \N__5054\,
            I => \N__4878\
        );

    \I__873\ : InMux
    port map (
            O => \N__5053\,
            I => \N__4878\
        );

    \I__872\ : InMux
    port map (
            O => \N__5052\,
            I => \N__4878\
        );

    \I__871\ : InMux
    port map (
            O => \N__5051\,
            I => \N__4878\
        );

    \I__870\ : InMux
    port map (
            O => \N__5050\,
            I => \N__4878\
        );

    \I__869\ : InMux
    port map (
            O => \N__5049\,
            I => \N__4878\
        );

    \I__868\ : InMux
    port map (
            O => \N__5048\,
            I => \N__4875\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__5045\,
            I => \N__4872\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5040\,
            I => \N__4867\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__5037\,
            I => \N__4867\
        );

    \I__864\ : InMux
    port map (
            O => \N__5036\,
            I => \N__4862\
        );

    \I__863\ : InMux
    port map (
            O => \N__5035\,
            I => \N__4862\
        );

    \I__862\ : InMux
    port map (
            O => \N__5034\,
            I => \N__4857\
        );

    \I__861\ : InMux
    port map (
            O => \N__5033\,
            I => \N__4854\
        );

    \I__860\ : Span4Mux_v
    port map (
            O => \N__5030\,
            I => \N__4849\
        );

    \I__859\ : Span4Mux_v
    port map (
            O => \N__5025\,
            I => \N__4849\
        );

    \I__858\ : Span4Mux_v
    port map (
            O => \N__5022\,
            I => \N__4844\
        );

    \I__857\ : Span4Mux_h
    port map (
            O => \N__5017\,
            I => \N__4844\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__5012\,
            I => \N__4841\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4999\,
            I => \N__4836\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__4986\,
            I => \N__4836\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4971\,
            I => \N__4833\
        );

    \I__852\ : Span4Mux_h
    port map (
            O => \N__4966\,
            I => \N__4822\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__4949\,
            I => \N__4822\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4932\,
            I => \N__4822\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__4915\,
            I => \N__4822\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4898\,
            I => \N__4822\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4895\,
            I => \N__4815\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4878\,
            I => \N__4815\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4875\,
            I => \N__4815\
        );

    \I__844\ : Span4Mux_v
    port map (
            O => \N__4872\,
            I => \N__4808\
        );

    \I__843\ : Span4Mux_h
    port map (
            O => \N__4867\,
            I => \N__4808\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4862\,
            I => \N__4808\
        );

    \I__841\ : InMux
    port map (
            O => \N__4861\,
            I => \N__4803\
        );

    \I__840\ : InMux
    port map (
            O => \N__4860\,
            I => \N__4803\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4857\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__4854\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__837\ : Odrv4
    port map (
            O => \N__4849\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__836\ : Odrv4
    port map (
            O => \N__4844\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__835\ : Odrv12
    port map (
            O => \N__4841\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__834\ : Odrv4
    port map (
            O => \N__4836\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__833\ : Odrv4
    port map (
            O => \N__4833\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__832\ : Odrv4
    port map (
            O => \N__4822\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__831\ : Odrv12
    port map (
            O => \N__4815\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__830\ : Odrv4
    port map (
            O => \N__4808\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__4803\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__828\ : CascadeMux
    port map (
            O => \N__4780\,
            I => \N__4777\
        );

    \I__827\ : InMux
    port map (
            O => \N__4777\,
            I => \N__4769\
        );

    \I__826\ : InMux
    port map (
            O => \N__4776\,
            I => \N__4739\
        );

    \I__825\ : InMux
    port map (
            O => \N__4775\,
            I => \N__4739\
        );

    \I__824\ : InMux
    port map (
            O => \N__4774\,
            I => \N__4739\
        );

    \I__823\ : InMux
    port map (
            O => \N__4773\,
            I => \N__4739\
        );

    \I__822\ : InMux
    port map (
            O => \N__4772\,
            I => \N__4736\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4769\,
            I => \N__4733\
        );

    \I__820\ : InMux
    port map (
            O => \N__4768\,
            I => \N__4730\
        );

    \I__819\ : InMux
    port map (
            O => \N__4767\,
            I => \N__4724\
        );

    \I__818\ : InMux
    port map (
            O => \N__4766\,
            I => \N__4724\
        );

    \I__817\ : InMux
    port map (
            O => \N__4765\,
            I => \N__4715\
        );

    \I__816\ : InMux
    port map (
            O => \N__4764\,
            I => \N__4715\
        );

    \I__815\ : InMux
    port map (
            O => \N__4763\,
            I => \N__4715\
        );

    \I__814\ : InMux
    port map (
            O => \N__4762\,
            I => \N__4715\
        );

    \I__813\ : InMux
    port map (
            O => \N__4761\,
            I => \N__4710\
        );

    \I__812\ : InMux
    port map (
            O => \N__4760\,
            I => \N__4710\
        );

    \I__811\ : InMux
    port map (
            O => \N__4759\,
            I => \N__4699\
        );

    \I__810\ : InMux
    port map (
            O => \N__4758\,
            I => \N__4699\
        );

    \I__809\ : InMux
    port map (
            O => \N__4757\,
            I => \N__4699\
        );

    \I__808\ : InMux
    port map (
            O => \N__4756\,
            I => \N__4699\
        );

    \I__807\ : InMux
    port map (
            O => \N__4755\,
            I => \N__4699\
        );

    \I__806\ : InMux
    port map (
            O => \N__4754\,
            I => \N__4684\
        );

    \I__805\ : InMux
    port map (
            O => \N__4753\,
            I => \N__4684\
        );

    \I__804\ : InMux
    port map (
            O => \N__4752\,
            I => \N__4684\
        );

    \I__803\ : InMux
    port map (
            O => \N__4751\,
            I => \N__4684\
        );

    \I__802\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4684\
        );

    \I__801\ : InMux
    port map (
            O => \N__4749\,
            I => \N__4684\
        );

    \I__800\ : InMux
    port map (
            O => \N__4748\,
            I => \N__4684\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4739\,
            I => \N__4681\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4736\,
            I => \N__4678\
        );

    \I__797\ : Span4Mux_v
    port map (
            O => \N__4733\,
            I => \N__4673\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__4730\,
            I => \N__4673\
        );

    \I__795\ : InMux
    port map (
            O => \N__4729\,
            I => \N__4670\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__4724\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_0\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__4715\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_0\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__4710\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_0\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__4699\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_0\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4684\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_0\
        );

    \I__789\ : Odrv4
    port map (
            O => \N__4681\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_0\
        );

    \I__788\ : Odrv12
    port map (
            O => \N__4678\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_0\
        );

    \I__787\ : Odrv4
    port map (
            O => \N__4673\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_0\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__4670\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_0\
        );

    \I__785\ : InMux
    port map (
            O => \N__4651\,
            I => \N__4648\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__4648\,
            I => \N__4617\
        );

    \I__783\ : ClkMux
    port map (
            O => \N__4647\,
            I => \N__4558\
        );

    \I__782\ : ClkMux
    port map (
            O => \N__4646\,
            I => \N__4558\
        );

    \I__781\ : ClkMux
    port map (
            O => \N__4645\,
            I => \N__4558\
        );

    \I__780\ : ClkMux
    port map (
            O => \N__4644\,
            I => \N__4558\
        );

    \I__779\ : ClkMux
    port map (
            O => \N__4643\,
            I => \N__4558\
        );

    \I__778\ : ClkMux
    port map (
            O => \N__4642\,
            I => \N__4558\
        );

    \I__777\ : ClkMux
    port map (
            O => \N__4641\,
            I => \N__4558\
        );

    \I__776\ : ClkMux
    port map (
            O => \N__4640\,
            I => \N__4558\
        );

    \I__775\ : ClkMux
    port map (
            O => \N__4639\,
            I => \N__4558\
        );

    \I__774\ : ClkMux
    port map (
            O => \N__4638\,
            I => \N__4558\
        );

    \I__773\ : ClkMux
    port map (
            O => \N__4637\,
            I => \N__4558\
        );

    \I__772\ : ClkMux
    port map (
            O => \N__4636\,
            I => \N__4558\
        );

    \I__771\ : ClkMux
    port map (
            O => \N__4635\,
            I => \N__4558\
        );

    \I__770\ : ClkMux
    port map (
            O => \N__4634\,
            I => \N__4558\
        );

    \I__769\ : ClkMux
    port map (
            O => \N__4633\,
            I => \N__4558\
        );

    \I__768\ : ClkMux
    port map (
            O => \N__4632\,
            I => \N__4558\
        );

    \I__767\ : ClkMux
    port map (
            O => \N__4631\,
            I => \N__4558\
        );

    \I__766\ : ClkMux
    port map (
            O => \N__4630\,
            I => \N__4558\
        );

    \I__765\ : ClkMux
    port map (
            O => \N__4629\,
            I => \N__4558\
        );

    \I__764\ : ClkMux
    port map (
            O => \N__4628\,
            I => \N__4558\
        );

    \I__763\ : ClkMux
    port map (
            O => \N__4627\,
            I => \N__4558\
        );

    \I__762\ : ClkMux
    port map (
            O => \N__4626\,
            I => \N__4558\
        );

    \I__761\ : ClkMux
    port map (
            O => \N__4625\,
            I => \N__4558\
        );

    \I__760\ : ClkMux
    port map (
            O => \N__4624\,
            I => \N__4558\
        );

    \I__759\ : ClkMux
    port map (
            O => \N__4623\,
            I => \N__4558\
        );

    \I__758\ : ClkMux
    port map (
            O => \N__4622\,
            I => \N__4558\
        );

    \I__757\ : ClkMux
    port map (
            O => \N__4621\,
            I => \N__4558\
        );

    \I__756\ : ClkMux
    port map (
            O => \N__4620\,
            I => \N__4558\
        );

    \I__755\ : Glb2LocalMux
    port map (
            O => \N__4617\,
            I => \N__4558\
        );

    \I__754\ : GlobalMux
    port map (
            O => \N__4558\,
            I => \N__4555\
        );

    \I__753\ : gio2CtrlBuf
    port map (
            O => \N__4555\,
            I => \CLK_c_g\
        );

    \I__752\ : InMux
    port map (
            O => \N__4552\,
            I => \N__4546\
        );

    \I__751\ : InMux
    port map (
            O => \N__4551\,
            I => \N__4546\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__4546\,
            I => \fsm_ctrl_inst1.toggle_clk_uCZ0Z1\
        );

    \I__749\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4540\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4540\,
            I => \N__4537\
        );

    \I__747\ : Odrv4
    port map (
            O => \N__4537\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_87\
        );

    \I__746\ : InMux
    port map (
            O => \N__4534\,
            I => \N__4531\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__4531\,
            I => \N__4528\
        );

    \I__744\ : Span4Mux_v
    port map (
            O => \N__4528\,
            I => \N__4524\
        );

    \I__743\ : InMux
    port map (
            O => \N__4527\,
            I => \N__4521\
        );

    \I__742\ : Odrv4
    port map (
            O => \N__4524\,
            I => \MOSI\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__4521\,
            I => \MOSI\
        );

    \I__740\ : InMux
    port map (
            O => \N__4516\,
            I => \N__4513\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__4513\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_85\
        );

    \I__738\ : InMux
    port map (
            O => \N__4510\,
            I => \N__4507\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__4507\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_86\
        );

    \I__736\ : InMux
    port map (
            O => \N__4504\,
            I => \N__4501\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__4501\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_0\
        );

    \I__734\ : InMux
    port map (
            O => \N__4498\,
            I => \N__4495\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4495\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_3\
        );

    \I__732\ : InMux
    port map (
            O => \N__4492\,
            I => \N__4489\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4489\,
            I => \N__4486\
        );

    \I__730\ : Odrv4
    port map (
            O => \N__4486\,
            I => \fsm_ctrl_inst1.current_state_ns_0_i_0_1_0\
        );

    \I__729\ : CascadeMux
    port map (
            O => \N__4483\,
            I => \N__4480\
        );

    \I__728\ : InMux
    port map (
            O => \N__4480\,
            I => \N__4477\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__4477\,
            I => \N__4474\
        );

    \I__726\ : Odrv4
    port map (
            O => \N__4474\,
            I => \fsm_ctrl_inst1.N_122_2\
        );

    \I__725\ : CascadeMux
    port map (
            O => \N__4471\,
            I => \N__4468\
        );

    \I__724\ : InMux
    port map (
            O => \N__4468\,
            I => \N__4464\
        );

    \I__723\ : InMux
    port map (
            O => \N__4467\,
            I => \N__4461\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4464\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_0\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__4461\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_0\
        );

    \I__720\ : InMux
    port map (
            O => \N__4456\,
            I => \bfn_7_25_0_\
        );

    \I__719\ : InMux
    port map (
            O => \N__4453\,
            I => \N__4448\
        );

    \I__718\ : InMux
    port map (
            O => \N__4452\,
            I => \N__4445\
        );

    \I__717\ : InMux
    port map (
            O => \N__4451\,
            I => \N__4442\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__4448\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_1\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__4445\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_1\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__4442\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_1\
        );

    \I__713\ : InMux
    port map (
            O => \N__4435\,
            I => \fsm_ctrl_inst1.counter_idle_cry_0\
        );

    \I__712\ : InMux
    port map (
            O => \N__4432\,
            I => \N__4427\
        );

    \I__711\ : InMux
    port map (
            O => \N__4431\,
            I => \N__4424\
        );

    \I__710\ : InMux
    port map (
            O => \N__4430\,
            I => \N__4421\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__4427\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_2\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__4424\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_2\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__4421\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_2\
        );

    \I__706\ : InMux
    port map (
            O => \N__4414\,
            I => \fsm_ctrl_inst1.counter_idle_cry_1\
        );

    \I__705\ : InMux
    port map (
            O => \N__4411\,
            I => \N__4406\
        );

    \I__704\ : InMux
    port map (
            O => \N__4410\,
            I => \N__4403\
        );

    \I__703\ : InMux
    port map (
            O => \N__4409\,
            I => \N__4400\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__4406\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_3\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__4403\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_3\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__4400\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_3\
        );

    \I__699\ : InMux
    port map (
            O => \N__4393\,
            I => \fsm_ctrl_inst1.counter_idle_cry_2\
        );

    \I__698\ : InMux
    port map (
            O => \N__4390\,
            I => \N__4381\
        );

    \I__697\ : InMux
    port map (
            O => \N__4389\,
            I => \N__4381\
        );

    \I__696\ : InMux
    port map (
            O => \N__4388\,
            I => \N__4374\
        );

    \I__695\ : InMux
    port map (
            O => \N__4387\,
            I => \N__4374\
        );

    \I__694\ : InMux
    port map (
            O => \N__4386\,
            I => \N__4374\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__4381\,
            I => \fsm_ctrl_inst1.current_state_23_d_i\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__4374\,
            I => \fsm_ctrl_inst1.current_state_23_d_i\
        );

    \I__691\ : InMux
    port map (
            O => \N__4369\,
            I => \fsm_ctrl_inst1.counter_idle_cry_3\
        );

    \I__690\ : CascadeMux
    port map (
            O => \N__4366\,
            I => \N__4361\
        );

    \I__689\ : InMux
    port map (
            O => \N__4365\,
            I => \N__4358\
        );

    \I__688\ : InMux
    port map (
            O => \N__4364\,
            I => \N__4355\
        );

    \I__687\ : InMux
    port map (
            O => \N__4361\,
            I => \N__4352\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4358\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_4\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4355\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_4\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__4352\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_4\
        );

    \I__683\ : CEMux
    port map (
            O => \N__4345\,
            I => \N__4342\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__4342\,
            I => \fsm_ctrl_inst1.counter_idlee_0_i\
        );

    \I__681\ : InMux
    port map (
            O => \N__4339\,
            I => \N__4336\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__4336\,
            I => \fsm_ctrl_inst1.toggle_clk_uC3Z0Z_0\
        );

    \I__679\ : InMux
    port map (
            O => \N__4333\,
            I => \N__4330\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__4330\,
            I => \N__4327\
        );

    \I__677\ : Odrv4
    port map (
            O => \N__4327\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_15\
        );

    \I__676\ : CascadeMux
    port map (
            O => \N__4324\,
            I => \N__4321\
        );

    \I__675\ : InMux
    port map (
            O => \N__4321\,
            I => \N__4318\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__4318\,
            I => \N__4315\
        );

    \I__673\ : Odrv4
    port map (
            O => \N__4315\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_87\
        );

    \I__672\ : InMux
    port map (
            O => \N__4312\,
            I => \N__4306\
        );

    \I__671\ : InMux
    port map (
            O => \N__4311\,
            I => \N__4306\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__4306\,
            I => \fsm_ctrl_inst1.N_119_0\
        );

    \I__669\ : CascadeMux
    port map (
            O => \N__4303\,
            I => \fsm_ctrl_inst1.N_105_cascade_\
        );

    \I__668\ : CascadeMux
    port map (
            O => \N__4300\,
            I => \N__4296\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__4299\,
            I => \N__4293\
        );

    \I__666\ : InMux
    port map (
            O => \N__4296\,
            I => \N__4288\
        );

    \I__665\ : InMux
    port map (
            O => \N__4293\,
            I => \N__4288\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__4288\,
            I => \fsm_ctrl_inst1.counter_dinZ0Z_3\
        );

    \I__663\ : CascadeMux
    port map (
            O => \N__4285\,
            I => \N__4282\
        );

    \I__662\ : InMux
    port map (
            O => \N__4282\,
            I => \N__4273\
        );

    \I__661\ : InMux
    port map (
            O => \N__4281\,
            I => \N__4273\
        );

    \I__660\ : InMux
    port map (
            O => \N__4280\,
            I => \N__4273\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__4273\,
            I => \fsm_ctrl_inst1.counter_dinZ0Z_2\
        );

    \I__658\ : InMux
    port map (
            O => \N__4270\,
            I => \N__4255\
        );

    \I__657\ : InMux
    port map (
            O => \N__4269\,
            I => \N__4255\
        );

    \I__656\ : InMux
    port map (
            O => \N__4268\,
            I => \N__4255\
        );

    \I__655\ : InMux
    port map (
            O => \N__4267\,
            I => \N__4255\
        );

    \I__654\ : InMux
    port map (
            O => \N__4266\,
            I => \N__4255\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__4255\,
            I => \fsm_ctrl_inst1.counter_dinZ0Z_0\
        );

    \I__652\ : CascadeMux
    port map (
            O => \N__4252\,
            I => \N__4248\
        );

    \I__651\ : InMux
    port map (
            O => \N__4251\,
            I => \N__4237\
        );

    \I__650\ : InMux
    port map (
            O => \N__4248\,
            I => \N__4237\
        );

    \I__649\ : InMux
    port map (
            O => \N__4247\,
            I => \N__4237\
        );

    \I__648\ : InMux
    port map (
            O => \N__4246\,
            I => \N__4237\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__4237\,
            I => \fsm_ctrl_inst1.counter_dinZ0Z_1\
        );

    \I__646\ : InMux
    port map (
            O => \N__4234\,
            I => \N__4231\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4231\,
            I => \N__4227\
        );

    \I__644\ : InMux
    port map (
            O => \N__4230\,
            I => \N__4224\
        );

    \I__643\ : Span4Mux_v
    port map (
            O => \N__4227\,
            I => \N__4218\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__4224\,
            I => \N__4218\
        );

    \I__641\ : InMux
    port map (
            O => \N__4223\,
            I => \N__4215\
        );

    \I__640\ : Odrv4
    port map (
            O => \N__4218\,
            I => \SEL_REG\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4215\,
            I => \SEL_REG\
        );

    \I__638\ : InMux
    port map (
            O => \N__4210\,
            I => \N__4207\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4207\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_15\
        );

    \I__636\ : IoInMux
    port map (
            O => \N__4204\,
            I => \N__4201\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__4201\,
            I => \N__4198\
        );

    \I__634\ : IoSpan4Mux
    port map (
            O => \N__4198\,
            I => \N__4195\
        );

    \I__633\ : Span4Mux_s3_h
    port map (
            O => \N__4195\,
            I => \N__4192\
        );

    \I__632\ : Span4Mux_v
    port map (
            O => \N__4192\,
            I => \N__4189\
        );

    \I__631\ : Sp12to4
    port map (
            O => \N__4189\,
            I => \N__4186\
        );

    \I__630\ : Span12Mux_v
    port map (
            O => \N__4186\,
            I => \N__4183\
        );

    \I__629\ : Odrv12
    port map (
            O => \N__4183\,
            I => \SDO_signal_out_c\
        );

    \I__628\ : InMux
    port map (
            O => \N__4180\,
            I => \N__4177\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__4177\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_36\
        );

    \I__626\ : InMux
    port map (
            O => \N__4174\,
            I => \N__4171\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__4171\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_37\
        );

    \I__624\ : InMux
    port map (
            O => \N__4168\,
            I => \N__4165\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__4165\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_50\
        );

    \I__622\ : InMux
    port map (
            O => \N__4162\,
            I => \N__4159\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__4159\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_51\
        );

    \I__620\ : InMux
    port map (
            O => \N__4156\,
            I => \N__4153\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__4153\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_38\
        );

    \I__618\ : InMux
    port map (
            O => \N__4150\,
            I => \N__4147\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__4147\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_39\
        );

    \I__616\ : InMux
    port map (
            O => \N__4144\,
            I => \N__4141\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__4141\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_86\
        );

    \I__614\ : InMux
    port map (
            O => \N__4138\,
            I => \N__4135\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__4135\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_17\
        );

    \I__612\ : InMux
    port map (
            O => \N__4132\,
            I => \N__4129\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__4129\,
            I => \N__4126\
        );

    \I__610\ : Odrv4
    port map (
            O => \N__4126\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_18\
        );

    \I__609\ : InMux
    port map (
            O => \N__4123\,
            I => \N__4120\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__4120\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_42\
        );

    \I__607\ : InMux
    port map (
            O => \N__4117\,
            I => \N__4114\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__4114\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_40\
        );

    \I__605\ : InMux
    port map (
            O => \N__4111\,
            I => \N__4108\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__4108\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_41\
        );

    \I__603\ : CEMux
    port map (
            O => \N__4105\,
            I => \N__4045\
        );

    \I__602\ : CEMux
    port map (
            O => \N__4104\,
            I => \N__4045\
        );

    \I__601\ : CEMux
    port map (
            O => \N__4103\,
            I => \N__4045\
        );

    \I__600\ : CEMux
    port map (
            O => \N__4102\,
            I => \N__4045\
        );

    \I__599\ : CEMux
    port map (
            O => \N__4101\,
            I => \N__4045\
        );

    \I__598\ : CEMux
    port map (
            O => \N__4100\,
            I => \N__4045\
        );

    \I__597\ : CEMux
    port map (
            O => \N__4099\,
            I => \N__4045\
        );

    \I__596\ : CEMux
    port map (
            O => \N__4098\,
            I => \N__4045\
        );

    \I__595\ : CEMux
    port map (
            O => \N__4097\,
            I => \N__4045\
        );

    \I__594\ : CEMux
    port map (
            O => \N__4096\,
            I => \N__4045\
        );

    \I__593\ : CEMux
    port map (
            O => \N__4095\,
            I => \N__4045\
        );

    \I__592\ : CEMux
    port map (
            O => \N__4094\,
            I => \N__4045\
        );

    \I__591\ : CEMux
    port map (
            O => \N__4093\,
            I => \N__4045\
        );

    \I__590\ : CEMux
    port map (
            O => \N__4092\,
            I => \N__4045\
        );

    \I__589\ : CEMux
    port map (
            O => \N__4091\,
            I => \N__4045\
        );

    \I__588\ : CEMux
    port map (
            O => \N__4090\,
            I => \N__4045\
        );

    \I__587\ : CEMux
    port map (
            O => \N__4089\,
            I => \N__4045\
        );

    \I__586\ : CEMux
    port map (
            O => \N__4088\,
            I => \N__4045\
        );

    \I__585\ : CEMux
    port map (
            O => \N__4087\,
            I => \N__4045\
        );

    \I__584\ : CEMux
    port map (
            O => \N__4086\,
            I => \N__4045\
        );

    \I__583\ : GlobalMux
    port map (
            O => \N__4045\,
            I => \N__4042\
        );

    \I__582\ : gio2CtrlBuf
    port map (
            O => \N__4042\,
            I => \fsm_ctrl_inst1.current_state_i_g_0\
        );

    \I__581\ : IoInMux
    port map (
            O => \N__4039\,
            I => \N__4036\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__4036\,
            I => \N__4033\
        );

    \I__579\ : Span4Mux_s3_h
    port map (
            O => \N__4033\,
            I => \N__4030\
        );

    \I__578\ : Span4Mux_v
    port map (
            O => \N__4030\,
            I => \N__4027\
        );

    \I__577\ : Odrv4
    port map (
            O => \N__4027\,
            I => \fsm_ctrl_inst1.current_state_i_0\
        );

    \I__576\ : CascadeMux
    port map (
            O => \N__4024\,
            I => \N__4019\
        );

    \I__575\ : InMux
    port map (
            O => \N__4023\,
            I => \N__4014\
        );

    \I__574\ : InMux
    port map (
            O => \N__4022\,
            I => \N__4014\
        );

    \I__573\ : InMux
    port map (
            O => \N__4019\,
            I => \N__4011\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4014\,
            I => \toggle_clk_uC4_0\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4011\,
            I => \toggle_clk_uC4_0\
        );

    \I__570\ : InMux
    port map (
            O => \N__4006\,
            I => \N__4002\
        );

    \I__569\ : InMux
    port map (
            O => \N__4005\,
            I => \N__3999\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__4002\,
            I => \fsm_ctrl_inst1_CLK_uC_1_i\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__3999\,
            I => \fsm_ctrl_inst1_CLK_uC_1_i\
        );

    \I__566\ : IoInMux
    port map (
            O => \N__3994\,
            I => \N__3991\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__3991\,
            I => \N__3988\
        );

    \I__564\ : Span4Mux_s3_v
    port map (
            O => \N__3988\,
            I => \N__3985\
        );

    \I__563\ : Span4Mux_v
    port map (
            O => \N__3985\,
            I => \N__3982\
        );

    \I__562\ : Sp12to4
    port map (
            O => \N__3982\,
            I => \N__3979\
        );

    \I__561\ : Odrv12
    port map (
            O => \N__3979\,
            I => \STATSR_cnv_0\
        );

    \I__560\ : CascadeMux
    port map (
            O => \N__3976\,
            I => \fsm_ctrl_inst1.counter_idlelde_0_a3_0_cascade_\
        );

    \I__559\ : InMux
    port map (
            O => \N__3973\,
            I => \N__3970\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__3970\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_78\
        );

    \I__557\ : InMux
    port map (
            O => \N__3967\,
            I => \N__3964\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__3964\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_79\
        );

    \I__555\ : InMux
    port map (
            O => \N__3961\,
            I => \N__3958\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3958\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_52\
        );

    \I__553\ : InMux
    port map (
            O => \N__3955\,
            I => \N__3952\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3952\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_35\
        );

    \I__551\ : InMux
    port map (
            O => \N__3949\,
            I => \N__3946\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__3946\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_49\
        );

    \I__549\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3940\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3940\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_0\
        );

    \I__547\ : InMux
    port map (
            O => \N__3937\,
            I => \N__3934\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3934\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_1\
        );

    \I__545\ : InMux
    port map (
            O => \N__3931\,
            I => \N__3928\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3928\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_9\
        );

    \I__543\ : InMux
    port map (
            O => \N__3925\,
            I => \N__3922\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3922\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_10\
        );

    \I__541\ : InMux
    port map (
            O => \N__3919\,
            I => \N__3916\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__3916\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_11\
        );

    \I__539\ : InMux
    port map (
            O => \N__3913\,
            I => \N__3910\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3910\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_12\
        );

    \I__537\ : InMux
    port map (
            O => \N__3907\,
            I => \N__3904\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3904\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_13\
        );

    \I__535\ : InMux
    port map (
            O => \N__3901\,
            I => \N__3898\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3898\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_14\
        );

    \I__533\ : CEMux
    port map (
            O => \N__3895\,
            I => \N__3891\
        );

    \I__532\ : CEMux
    port map (
            O => \N__3894\,
            I => \N__3888\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3891\,
            I => \N__3885\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3888\,
            I => \N__3882\
        );

    \I__529\ : Span4Mux_v
    port map (
            O => \N__3885\,
            I => \N__3879\
        );

    \I__528\ : Odrv12
    port map (
            O => \N__3882\,
            I => \config_register_latched_dec_inst1.DYNSR_cnvZ0Z_0\
        );

    \I__527\ : Odrv4
    port map (
            O => \N__3879\,
            I => \config_register_latched_dec_inst1.DYNSR_cnvZ0Z_0\
        );

    \I__526\ : InMux
    port map (
            O => \N__3874\,
            I => \fsm_ctrl_inst1.counter_stat_cry_2\
        );

    \I__525\ : InMux
    port map (
            O => \N__3871\,
            I => \fsm_ctrl_inst1.counter_stat_cry_3\
        );

    \I__524\ : InMux
    port map (
            O => \N__3868\,
            I => \fsm_ctrl_inst1.counter_stat_cry_4\
        );

    \I__523\ : CEMux
    port map (
            O => \N__3865\,
            I => \N__3857\
        );

    \I__522\ : CEMux
    port map (
            O => \N__3864\,
            I => \N__3854\
        );

    \I__521\ : InMux
    port map (
            O => \N__3863\,
            I => \N__3847\
        );

    \I__520\ : InMux
    port map (
            O => \N__3862\,
            I => \N__3847\
        );

    \I__519\ : InMux
    port map (
            O => \N__3861\,
            I => \N__3847\
        );

    \I__518\ : CEMux
    port map (
            O => \N__3860\,
            I => \N__3840\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3857\,
            I => \N__3837\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3854\,
            I => \N__3834\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3847\,
            I => \N__3831\
        );

    \I__514\ : InMux
    port map (
            O => \N__3846\,
            I => \N__3822\
        );

    \I__513\ : InMux
    port map (
            O => \N__3845\,
            I => \N__3822\
        );

    \I__512\ : InMux
    port map (
            O => \N__3844\,
            I => \N__3822\
        );

    \I__511\ : InMux
    port map (
            O => \N__3843\,
            I => \N__3822\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__3840\,
            I => \N__3819\
        );

    \I__509\ : Span4Mux_v
    port map (
            O => \N__3837\,
            I => \N__3816\
        );

    \I__508\ : Span4Mux_h
    port map (
            O => \N__3834\,
            I => \N__3813\
        );

    \I__507\ : Odrv4
    port map (
            O => \N__3831\,
            I => \fsm_ctrl_inst1.current_state_i_1\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3822\,
            I => \fsm_ctrl_inst1.current_state_i_1\
        );

    \I__505\ : Odrv12
    port map (
            O => \N__3819\,
            I => \fsm_ctrl_inst1.current_state_i_1\
        );

    \I__504\ : Odrv4
    port map (
            O => \N__3816\,
            I => \fsm_ctrl_inst1.current_state_i_1\
        );

    \I__503\ : Odrv4
    port map (
            O => \N__3813\,
            I => \fsm_ctrl_inst1.current_state_i_1\
        );

    \I__502\ : InMux
    port map (
            O => \N__3802\,
            I => \fsm_ctrl_inst1.counter_stat_cry_5\
        );

    \I__501\ : CEMux
    port map (
            O => \N__3799\,
            I => \N__3796\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3796\,
            I => \fsm_ctrl_inst1.counter_state_0_i\
        );

    \I__499\ : InMux
    port map (
            O => \N__3793\,
            I => \N__3788\
        );

    \I__498\ : InMux
    port map (
            O => \N__3792\,
            I => \N__3785\
        );

    \I__497\ : InMux
    port map (
            O => \N__3791\,
            I => \N__3782\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__3788\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_3\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__3785\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_3\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3782\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_3\
        );

    \I__493\ : InMux
    port map (
            O => \N__3775\,
            I => \N__3771\
        );

    \I__492\ : InMux
    port map (
            O => \N__3774\,
            I => \N__3768\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3771\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_1\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3768\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_1\
        );

    \I__489\ : CascadeMux
    port map (
            O => \N__3763\,
            I => \N__3759\
        );

    \I__488\ : InMux
    port map (
            O => \N__3762\,
            I => \N__3755\
        );

    \I__487\ : InMux
    port map (
            O => \N__3759\,
            I => \N__3752\
        );

    \I__486\ : InMux
    port map (
            O => \N__3758\,
            I => \N__3749\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3755\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_6\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3752\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_6\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__3749\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_6\
        );

    \I__482\ : InMux
    port map (
            O => \N__3742\,
            I => \N__3738\
        );

    \I__481\ : InMux
    port map (
            O => \N__3741\,
            I => \N__3735\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3738\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_0\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__3735\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_0\
        );

    \I__478\ : InMux
    port map (
            O => \N__3730\,
            I => \N__3725\
        );

    \I__477\ : InMux
    port map (
            O => \N__3729\,
            I => \N__3722\
        );

    \I__476\ : InMux
    port map (
            O => \N__3728\,
            I => \N__3719\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__3725\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_5\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__3722\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_5\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3719\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_5\
        );

    \I__472\ : InMux
    port map (
            O => \N__3712\,
            I => \N__3708\
        );

    \I__471\ : InMux
    port map (
            O => \N__3711\,
            I => \N__3705\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3708\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_2\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3705\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_2\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__3700\,
            I => \fsm_ctrl_inst1.current_state_ns_i_a3_0_4_1_cascade_\
        );

    \I__467\ : InMux
    port map (
            O => \N__3697\,
            I => \N__3692\
        );

    \I__466\ : InMux
    port map (
            O => \N__3696\,
            I => \N__3689\
        );

    \I__465\ : InMux
    port map (
            O => \N__3695\,
            I => \N__3686\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3692\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_4\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__3689\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_4\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3686\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_4\
        );

    \I__461\ : CascadeMux
    port map (
            O => \N__3679\,
            I => \fsm_ctrl_inst1.current_state_ns_i_a3_0_5_1_cascade_\
        );

    \I__460\ : InMux
    port map (
            O => \N__3676\,
            I => \N__3673\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3673\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_15\
        );

    \I__458\ : InMux
    port map (
            O => \N__3670\,
            I => \N__3667\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3667\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_16\
        );

    \I__456\ : InMux
    port map (
            O => \N__3664\,
            I => \N__3661\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__3661\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_5\
        );

    \I__454\ : InMux
    port map (
            O => \N__3658\,
            I => \N__3655\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3655\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_6\
        );

    \I__452\ : InMux
    port map (
            O => \N__3652\,
            I => \N__3649\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__3649\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_45\
        );

    \I__450\ : InMux
    port map (
            O => \N__3646\,
            I => \N__3643\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__3643\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_46\
        );

    \I__448\ : InMux
    port map (
            O => \N__3640\,
            I => \N__3637\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__3637\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_43\
        );

    \I__446\ : InMux
    port map (
            O => \N__3634\,
            I => \N__3631\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__3631\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_44\
        );

    \I__444\ : InMux
    port map (
            O => \N__3628\,
            I => \bfn_6_21_0_\
        );

    \I__443\ : InMux
    port map (
            O => \N__3625\,
            I => \fsm_ctrl_inst1.counter_stat_cry_0\
        );

    \I__442\ : InMux
    port map (
            O => \N__3622\,
            I => \fsm_ctrl_inst1.counter_stat_cry_1\
        );

    \I__441\ : InMux
    port map (
            O => \N__3619\,
            I => \N__3616\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__3616\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_48\
        );

    \I__439\ : InMux
    port map (
            O => \N__3613\,
            I => \N__3610\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__3610\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_47\
        );

    \I__437\ : InMux
    port map (
            O => \N__3607\,
            I => \N__3604\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3604\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_59\
        );

    \I__435\ : InMux
    port map (
            O => \N__3601\,
            I => \N__3598\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__3598\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_60\
        );

    \I__433\ : InMux
    port map (
            O => \N__3595\,
            I => \N__3592\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__3592\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_85\
        );

    \I__431\ : InMux
    port map (
            O => \N__3589\,
            I => \N__3586\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__3586\,
            I => \N__3583\
        );

    \I__429\ : Odrv4
    port map (
            O => \N__3583\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_34\
        );

    \I__428\ : InMux
    port map (
            O => \N__3580\,
            I => \N__3577\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3577\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_80\
        );

    \I__426\ : InMux
    port map (
            O => \N__3574\,
            I => \N__3571\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__3571\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_3\
        );

    \I__424\ : InMux
    port map (
            O => \N__3568\,
            I => \N__3565\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__3565\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_4\
        );

    \I__422\ : InMux
    port map (
            O => \N__3562\,
            I => \N__3559\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3559\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_58\
        );

    \I__420\ : InMux
    port map (
            O => \N__3556\,
            I => \N__3553\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__3553\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_53\
        );

    \I__418\ : CascadeMux
    port map (
            O => \N__3550\,
            I => \N__3547\
        );

    \I__417\ : InMux
    port map (
            O => \N__3547\,
            I => \N__3544\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__3544\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_77\
        );

    \I__415\ : InMux
    port map (
            O => \N__3541\,
            I => \N__3538\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__3538\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_56\
        );

    \I__413\ : InMux
    port map (
            O => \N__3535\,
            I => \N__3532\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__3532\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_57\
        );

    \I__411\ : InMux
    port map (
            O => \N__3529\,
            I => \N__3526\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__3526\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_54\
        );

    \I__409\ : InMux
    port map (
            O => \N__3523\,
            I => \N__3520\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__3520\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_55\
        );

    \I__407\ : InMux
    port map (
            O => \N__3517\,
            I => \N__3514\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__3514\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_3\
        );

    \I__405\ : InMux
    port map (
            O => \N__3511\,
            I => \N__3508\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__3508\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_4\
        );

    \I__403\ : InMux
    port map (
            O => \N__3505\,
            I => \N__3502\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__3502\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_5\
        );

    \I__401\ : InMux
    port map (
            O => \N__3499\,
            I => \N__3496\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__3496\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_6\
        );

    \I__399\ : InMux
    port map (
            O => \N__3493\,
            I => \N__3490\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__3490\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_2\
        );

    \I__397\ : InMux
    port map (
            O => \N__3487\,
            I => \N__3484\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__3484\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_7\
        );

    \I__395\ : InMux
    port map (
            O => \N__3481\,
            I => \N__3478\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3478\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_8\
        );

    \I__393\ : InMux
    port map (
            O => \N__3475\,
            I => \N__3472\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__3472\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_76\
        );

    \I__391\ : InMux
    port map (
            O => \N__3469\,
            I => \N__3466\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3466\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_6\
        );

    \I__389\ : InMux
    port map (
            O => \N__3463\,
            I => \N__3460\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__3460\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_7\
        );

    \I__387\ : InMux
    port map (
            O => \N__3457\,
            I => \N__3454\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__3454\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_5\
        );

    \I__385\ : CascadeMux
    port map (
            O => \N__3451\,
            I => \fsm_ctrl_inst1.un1_counter_statlt5_0_cascade_\
        );

    \I__384\ : InMux
    port map (
            O => \N__3448\,
            I => \N__3445\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__3445\,
            I => \N__3442\
        );

    \I__382\ : Odrv4
    port map (
            O => \N__3442\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_4\
        );

    \I__381\ : InMux
    port map (
            O => \N__3439\,
            I => \N__3436\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__3436\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_2\
        );

    \I__379\ : InMux
    port map (
            O => \N__3433\,
            I => \N__3430\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__3430\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_3\
        );

    \I__377\ : InMux
    port map (
            O => \N__3427\,
            I => \N__3424\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__3424\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_0\
        );

    \I__375\ : InMux
    port map (
            O => \N__3421\,
            I => \N__3418\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__3418\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_1\
        );

    \I__373\ : InMux
    port map (
            O => \N__3415\,
            I => \N__3412\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__3412\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_62\
        );

    \I__371\ : InMux
    port map (
            O => \N__3409\,
            I => \N__3406\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__3406\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_2\
        );

    \I__369\ : InMux
    port map (
            O => \N__3403\,
            I => \N__3400\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__3400\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_8\
        );

    \I__367\ : InMux
    port map (
            O => \N__3397\,
            I => \N__3394\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__3394\,
            I => \N__3391\
        );

    \I__365\ : Odrv4
    port map (
            O => \N__3391\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_9\
        );

    \I__364\ : InMux
    port map (
            O => \N__3388\,
            I => \N__3385\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__3385\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_61\
        );

    \I__362\ : InMux
    port map (
            O => \N__3382\,
            I => \N__3379\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__3379\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_10\
        );

    \I__360\ : InMux
    port map (
            O => \N__3376\,
            I => \N__3373\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__3373\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_11\
        );

    \I__358\ : InMux
    port map (
            O => \N__3370\,
            I => \N__3367\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__3367\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_8\
        );

    \I__356\ : InMux
    port map (
            O => \N__3364\,
            I => \N__3361\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__3361\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_9\
        );

    \I__354\ : InMux
    port map (
            O => \N__3358\,
            I => \N__3355\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__3355\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_31\
        );

    \I__352\ : InMux
    port map (
            O => \N__3352\,
            I => \N__3349\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__3349\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_32\
        );

    \I__350\ : InMux
    port map (
            O => \N__3346\,
            I => \N__3343\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__3343\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_33\
        );

    \I__348\ : InMux
    port map (
            O => \N__3340\,
            I => \N__3337\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__3337\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_1\
        );

    \I__346\ : InMux
    port map (
            O => \N__3334\,
            I => \N__3331\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__3331\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_81\
        );

    \I__344\ : InMux
    port map (
            O => \N__3328\,
            I => \N__3325\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__3325\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_0\
        );

    \I__342\ : InMux
    port map (
            O => \N__3322\,
            I => \N__3319\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__3319\,
            I => \N__3316\
        );

    \I__340\ : Odrv4
    port map (
            O => \N__3316\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_19\
        );

    \I__339\ : InMux
    port map (
            O => \N__3313\,
            I => \N__3310\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__3310\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_7\
        );

    \I__337\ : InMux
    port map (
            O => \N__3307\,
            I => \N__3304\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__3304\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_14\
        );

    \I__335\ : InMux
    port map (
            O => \N__3301\,
            I => \N__3298\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__3298\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_12\
        );

    \I__333\ : InMux
    port map (
            O => \N__3295\,
            I => \N__3292\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__3292\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_13\
        );

    \I__331\ : InMux
    port map (
            O => \N__3289\,
            I => \N__3286\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__3286\,
            I => \N__3283\
        );

    \I__329\ : Odrv4
    port map (
            O => \N__3283\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_73\
        );

    \I__328\ : InMux
    port map (
            O => \N__3280\,
            I => \N__3277\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__3277\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_84\
        );

    \I__326\ : InMux
    port map (
            O => \N__3274\,
            I => \N__3271\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__3271\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_82\
        );

    \I__324\ : InMux
    port map (
            O => \N__3268\,
            I => \N__3265\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__3265\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_74\
        );

    \I__322\ : InMux
    port map (
            O => \N__3262\,
            I => \N__3259\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__3259\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_75\
        );

    \I__320\ : InMux
    port map (
            O => \N__3256\,
            I => \N__3253\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__3253\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_14\
        );

    \I__318\ : InMux
    port map (
            O => \N__3250\,
            I => \N__3247\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__3247\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_13\
        );

    \I__316\ : InMux
    port map (
            O => \N__3244\,
            I => \N__3241\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__3241\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_29\
        );

    \I__314\ : InMux
    port map (
            O => \N__3238\,
            I => \N__3235\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__3235\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_30\
        );

    \I__312\ : InMux
    port map (
            O => \N__3232\,
            I => \N__3229\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__3229\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_12\
        );

    \I__310\ : InMux
    port map (
            O => \N__3226\,
            I => \N__3223\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__3223\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_11\
        );

    \I__308\ : InMux
    port map (
            O => \N__3220\,
            I => \N__3217\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__3217\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_10\
        );

    \I__306\ : InMux
    port map (
            O => \N__3214\,
            I => \N__3211\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__3211\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_63\
        );

    \I__304\ : InMux
    port map (
            O => \N__3208\,
            I => \N__3205\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__3205\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_24\
        );

    \I__302\ : InMux
    port map (
            O => \N__3202\,
            I => \N__3199\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__3199\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_22\
        );

    \I__300\ : InMux
    port map (
            O => \N__3196\,
            I => \N__3193\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__3193\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_23\
        );

    \I__298\ : InMux
    port map (
            O => \N__3190\,
            I => \N__3187\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__3187\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_66\
        );

    \I__296\ : InMux
    port map (
            O => \N__3184\,
            I => \N__3181\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__3181\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_67\
        );

    \I__294\ : InMux
    port map (
            O => \N__3178\,
            I => \N__3175\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__3175\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_68\
        );

    \I__292\ : InMux
    port map (
            O => \N__3172\,
            I => \N__3169\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__3169\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_64\
        );

    \I__290\ : InMux
    port map (
            O => \N__3166\,
            I => \N__3163\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__3163\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_65\
        );

    \I__288\ : InMux
    port map (
            O => \N__3160\,
            I => \N__3157\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__3157\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_83\
        );

    \I__286\ : InMux
    port map (
            O => \N__3154\,
            I => \N__3151\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__3151\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_28\
        );

    \I__284\ : InMux
    port map (
            O => \N__3148\,
            I => \N__3145\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__3145\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_70\
        );

    \I__282\ : InMux
    port map (
            O => \N__3142\,
            I => \N__3139\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__3139\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_71\
        );

    \I__280\ : InMux
    port map (
            O => \N__3136\,
            I => \N__3133\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__3133\,
            I => \N__3130\
        );

    \I__278\ : Odrv4
    port map (
            O => \N__3130\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_20\
        );

    \I__277\ : InMux
    port map (
            O => \N__3127\,
            I => \N__3124\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__3124\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_26\
        );

    \I__275\ : InMux
    port map (
            O => \N__3121\,
            I => \N__3118\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__3118\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_27\
        );

    \I__273\ : InMux
    port map (
            O => \N__3115\,
            I => \N__3112\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__3112\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_69\
        );

    \I__271\ : InMux
    port map (
            O => \N__3109\,
            I => \N__3106\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__3106\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_25\
        );

    \I__269\ : InMux
    port map (
            O => \N__3103\,
            I => \N__3100\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__3100\,
            I => \RST_N_c\
        );

    \I__267\ : IoInMux
    port map (
            O => \N__3097\,
            I => \N__3094\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__3094\,
            I => \RST_N_c_i\
        );

    \I__265\ : InMux
    port map (
            O => \N__3091\,
            I => \N__3088\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__3088\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_21\
        );

    \I__263\ : InMux
    port map (
            O => \N__3085\,
            I => \N__3082\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__3082\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_72\
        );

    \IN_MUX_bfv_6_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_21_0_\
        );

    \IN_MUX_bfv_7_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_25_0_\
        );

    \fsm_ctrl_inst1.current_state_RNI1GR8_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4039\,
            GLOBALBUFFEROUTPUT => \fsm_ctrl_inst1.current_state_i_g_0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \RST_N_ibuf_RNIBJGC_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3097\,
            GLOBALBUFFEROUTPUT => \RST_N_c_i_g\
        );

    \N_224_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3994\,
            GLOBALBUFFEROUTPUT => \N_224_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \RST_N_ibuf_RNIBJGC_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3103\,
            lcout => \RST_N_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_22_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5118\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3091\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4636\,
            ce => \N__4093\,
            sr => \N__5761\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_21_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1011101110111011"
        )
    port map (
            in0 => \N__3136\,
            in1 => \N__5117\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4636\,
            ce => \N__4093\,
            sr => \N__5761\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_73_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3085\,
            in2 => \_gnd_net_\,
            in3 => \N__5171\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4647\,
            ce => \N__4086\,
            sr => \N__5754\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_72_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3142\,
            in2 => \_gnd_net_\,
            in3 => \N__5190\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4645\,
            ce => \N__4087\,
            sr => \N__5755\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_28_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3121\,
            in2 => \_gnd_net_\,
            in3 => \N__5188\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4645\,
            ce => \N__4087\,
            sr => \N__5755\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_29_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3154\,
            in2 => \_gnd_net_\,
            in3 => \N__5189\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4645\,
            ce => \N__4087\,
            sr => \N__5755\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_26_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3109\,
            in2 => \_gnd_net_\,
            in3 => \N__5177\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4641\,
            ce => \N__4090\,
            sr => \N__5757\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_70_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5179\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3115\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4641\,
            ce => \N__4090\,
            sr => \N__5757\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_71_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5180\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3148\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4641\,
            ce => \N__4090\,
            sr => \N__5757\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_20_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3322\,
            in2 => \_gnd_net_\,
            in3 => \N__5176\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4641\,
            ce => \N__4090\,
            sr => \N__5757\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_27_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5178\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3127\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4641\,
            ce => \N__4090\,
            sr => \N__5757\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_69_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5167\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3178\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4637\,
            ce => \N__4094\,
            sr => \N__5762\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_25_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3208\,
            in2 => \_gnd_net_\,
            in3 => \N__5166\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4637\,
            ce => \N__4094\,
            sr => \N__5762\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_64_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5100\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3214\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4631\,
            ce => \N__4098\,
            sr => \N__5766\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_24_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3196\,
            in2 => \_gnd_net_\,
            in3 => \N__5099\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4631\,
            ce => \N__4098\,
            sr => \N__5766\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_67_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5103\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3190\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4631\,
            ce => \N__4098\,
            sr => \N__5766\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_23_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3202\,
            in2 => \_gnd_net_\,
            in3 => \N__5098\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4631\,
            ce => \N__4098\,
            sr => \N__5766\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_66_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5102\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3166\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4631\,
            ce => \N__4098\,
            sr => \N__5766\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_68_LC_3_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5104\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3184\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4631\,
            ce => \N__4098\,
            sr => \N__5766\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_65_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3172\,
            in2 => \_gnd_net_\,
            in3 => \N__5101\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4631\,
            ce => \N__4098\,
            sr => \N__5766\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_83_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3274\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5169\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4646\,
            ce => \N__4088\,
            sr => \N__5756\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_84_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__5170\,
            in1 => \N__3160\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4646\,
            ce => \N__4088\,
            sr => \N__5756\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_34_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5187\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3346\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4642\,
            ce => \N__4091\,
            sr => \N__5758\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_14_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5185\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3250\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4642\,
            ce => \N__4091\,
            sr => \N__5758\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_31_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3238\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4642\,
            ce => \N__4091\,
            sr => \N__5758\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_13_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3232\,
            in2 => \_gnd_net_\,
            in3 => \N__5184\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4642\,
            ce => \N__4091\,
            sr => \N__5758\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_30_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__3244\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5175\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4638\,
            ce => \N__4095\,
            sr => \N__5763\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_12_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5174\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3226\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4638\,
            ce => \N__4095\,
            sr => \N__5763\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_11_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5173\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3220\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4638\,
            ce => \N__4095\,
            sr => \N__5763\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_10_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3397\,
            in2 => \_gnd_net_\,
            in3 => \N__5172\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4638\,
            ce => \N__4095\,
            sr => \N__5763\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_63_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3415\,
            in2 => \_gnd_net_\,
            in3 => \N__5165\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4632\,
            ce => \N__4099\,
            sr => \N__5767\
        );

    \fsm_ctrl_inst1.bit_sequence_din_14_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3295\,
            in2 => \_gnd_net_\,
            in3 => \N__4776\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4627\,
            ce => \N__3865\,
            sr => \N__5771\
        );

    \fsm_ctrl_inst1.bit_sequence_din_15_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4773\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3307\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4627\,
            ce => \N__3865\,
            sr => \N__5771\
        );

    \fsm_ctrl_inst1.bit_sequence_din_12_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3376\,
            in2 => \_gnd_net_\,
            in3 => \N__4774\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4627\,
            ce => \N__3865\,
            sr => \N__5771\
        );

    \fsm_ctrl_inst1.bit_sequence_din_13_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3301\,
            in2 => \_gnd_net_\,
            in3 => \N__4775\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4627\,
            ce => \N__3865\,
            sr => \N__5771\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_74_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3289\,
            in2 => \_gnd_net_\,
            in3 => \N__5181\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4643\,
            ce => \N__4092\,
            sr => \N__5759\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_76_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5182\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3262\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4643\,
            ce => \N__4092\,
            sr => \N__5759\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_85_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3280\,
            in2 => \_gnd_net_\,
            in3 => \N__5183\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4643\,
            ce => \N__4092\,
            sr => \N__5759\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_82_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5089\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3334\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4639\,
            ce => \N__4096\,
            sr => \N__5764\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_75_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3268\,
            in2 => \_gnd_net_\,
            in3 => \N__5087\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4639\,
            ce => \N__4096\,
            sr => \N__5764\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_15_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5082\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3256\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4639\,
            ce => \N__4096\,
            sr => \N__5764\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_32_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3358\,
            in2 => \_gnd_net_\,
            in3 => \N__5085\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4639\,
            ce => \N__4096\,
            sr => \N__5764\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_1_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__5083\,
            in1 => \N__3328\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4639\,
            ce => \N__4096\,
            sr => \N__5764\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_33_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3352\,
            in2 => \_gnd_net_\,
            in3 => \N__5086\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4639\,
            ce => \N__4096\,
            sr => \N__5764\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_2_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5084\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3340\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4639\,
            ce => \N__4096\,
            sr => \N__5764\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_81_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3580\,
            in2 => \_gnd_net_\,
            in3 => \N__5088\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4639\,
            ce => \N__4096\,
            sr => \N__5764\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_7_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5063\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3658\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4633\,
            ce => \N__4100\,
            sr => \N__5768\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_0_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5058\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4633\,
            ce => \N__4100\,
            sr => \N__5768\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_19_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5059\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4132\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4633\,
            ce => \N__4100\,
            sr => \N__5768\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_8_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3313\,
            in2 => \_gnd_net_\,
            in3 => \N__5064\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4633\,
            ce => \N__4100\,
            sr => \N__5768\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_62_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5062\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3388\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4633\,
            ce => \N__4100\,
            sr => \N__5768\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_3_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3409\,
            in2 => \_gnd_net_\,
            in3 => \N__5060\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4633\,
            ce => \N__4100\,
            sr => \N__5768\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_9_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5065\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3403\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4633\,
            ce => \N__4100\,
            sr => \N__5768\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_61_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3601\,
            in2 => \_gnd_net_\,
            in3 => \N__5061\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4633\,
            ce => \N__4100\,
            sr => \N__5768\
        );

    \fsm_ctrl_inst1.bit_sequence_din_6_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3457\,
            in2 => \_gnd_net_\,
            in3 => \N__4753\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4628\,
            ce => \N__3860\,
            sr => \N__5772\
        );

    \fsm_ctrl_inst1.bit_sequence_din_8_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4750\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3463\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4628\,
            ce => \N__3860\,
            sr => \N__5772\
        );

    \fsm_ctrl_inst1.bit_sequence_din_10_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3364\,
            in2 => \_gnd_net_\,
            in3 => \N__4751\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4628\,
            ce => \N__3860\,
            sr => \N__5772\
        );

    \fsm_ctrl_inst1.bit_sequence_din_11_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4748\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3382\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4628\,
            ce => \N__3860\,
            sr => \N__5772\
        );

    \fsm_ctrl_inst1.bit_sequence_din_9_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3370\,
            in2 => \_gnd_net_\,
            in3 => \N__4754\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4628\,
            ce => \N__3860\,
            sr => \N__5772\
        );

    \fsm_ctrl_inst1.bit_sequence_din_7_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4749\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3469\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4628\,
            ce => \N__3860\,
            sr => \N__5772\
        );

    \fsm_ctrl_inst1.bit_sequence_din_5_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3448\,
            in2 => \_gnd_net_\,
            in3 => \N__4752\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4628\,
            ce => \N__3860\,
            sr => \N__5772\
        );

    \fsm_ctrl_inst1.current_state_RNI2HR8_1_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4860\,
            lcout => \fsm_ctrl_inst1.current_state_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_stat_RNIPO4_3_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3695\,
            in2 => \_gnd_net_\,
            in3 => \N__3792\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.un1_counter_statlt5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_stat_RNIO659_6_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011111111111"
        )
    port map (
            in0 => \N__3730\,
            in1 => \N__4861\,
            in2 => \N__3451\,
            in3 => \N__3758\,
            lcout => \fsm_ctrl_inst1.counter_state_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.bit_sequence_din_4_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4757\,
            in2 => \_gnd_net_\,
            in3 => \N__3433\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4623\,
            ce => \N__3864\,
            sr => \N__5777\
        );

    \fsm_ctrl_inst1.bit_sequence_din_0_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4758\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4623\,
            ce => \N__3864\,
            sr => \N__5777\
        );

    \fsm_ctrl_inst1.bit_sequence_din_2_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4756\,
            in2 => \_gnd_net_\,
            in3 => \N__3421\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4623\,
            ce => \N__3864\,
            sr => \N__5777\
        );

    \fsm_ctrl_inst1.bit_sequence_din_3_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__4759\,
            in1 => \N__3439\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4623\,
            ce => \N__3864\,
            sr => \N__5777\
        );

    \fsm_ctrl_inst1.bit_sequence_din_1_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4755\,
            in2 => \_gnd_net_\,
            in3 => \N__3427\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4623\,
            ce => \N__3864\,
            sr => \N__5777\
        );

    \config_register_latched_dec_inst1.DYNSR_4_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3517\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5965\,
            ce => \N__3895\,
            sr => \N__5779\
        );

    \config_register_latched_dec_inst1.DYNSR_3_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3493\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5965\,
            ce => \N__3895\,
            sr => \N__5779\
        );

    \config_register_latched_dec_inst1.DYNSR_7_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3499\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5965\,
            ce => \N__3895\,
            sr => \N__5779\
        );

    \config_register_latched_dec_inst1.DYNSR_5_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3511\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5965\,
            ce => \N__3895\,
            sr => \N__5779\
        );

    \config_register_latched_dec_inst1.DYNSR_6_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3505\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5965\,
            ce => \N__3895\,
            sr => \N__5779\
        );

    \config_register_latched_dec_inst1.DYNSR_2_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3937\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5965\,
            ce => \N__3895\,
            sr => \N__5779\
        );

    \config_register_latched_dec_inst1.DYNSR_9_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3481\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5965\,
            ce => \N__3895\,
            sr => \N__5779\
        );

    \config_register_latched_dec_inst1.DYNSR_8_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3487\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5965\,
            ce => \N__3895\,
            sr => \N__5779\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_77_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__3475\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5057\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4644\,
            ce => \N__4089\,
            sr => \N__5760\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_59_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3562\,
            in2 => \_gnd_net_\,
            in3 => \N__5055\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4640\,
            ce => \N__4097\,
            sr => \N__5765\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_56_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5052\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3523\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4640\,
            ce => \N__4097\,
            sr => \N__5765\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_54_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3556\,
            in2 => \_gnd_net_\,
            in3 => \N__5050\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4640\,
            ce => \N__4097\,
            sr => \N__5765\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_58_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5054\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3535\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4640\,
            ce => \N__4097\,
            sr => \N__5765\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_53_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3961\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5049\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4640\,
            ce => \N__4097\,
            sr => \N__5765\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_78_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__5056\,
            in1 => \_gnd_net_\,
            in2 => \N__3550\,
            in3 => \_gnd_net_\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4640\,
            ce => \N__4097\,
            sr => \N__5765\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_57_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3541\,
            in2 => \_gnd_net_\,
            in3 => \N__5053\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4640\,
            ce => \N__4097\,
            sr => \N__5765\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_55_LC_6_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5051\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3529\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4640\,
            ce => \N__4097\,
            sr => \N__5765\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_5_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3568\,
            in2 => \_gnd_net_\,
            in3 => \N__5078\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4634\,
            ce => \N__4101\,
            sr => \N__5769\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_48_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5076\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3613\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4634\,
            ce => \N__4101\,
            sr => \N__5769\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_49_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3619\,
            in2 => \_gnd_net_\,
            in3 => \N__5077\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4634\,
            ce => \N__4101\,
            sr => \N__5769\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_47_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5075\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3646\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4634\,
            ce => \N__4101\,
            sr => \N__5769\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_60_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__3607\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5079\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4634\,
            ce => \N__4101\,
            sr => \N__5769\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_86_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5081\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3595\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4634\,
            ce => \N__4101\,
            sr => \N__5769\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_35_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3589\,
            in2 => \_gnd_net_\,
            in3 => \N__5074\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4634\,
            ce => \N__4101\,
            sr => \N__5769\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_80_LC_6_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5080\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3967\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4634\,
            ce => \N__4101\,
            sr => \N__5769\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_4_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3574\,
            in2 => \_gnd_net_\,
            in3 => \N__5072\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4629\,
            ce => \N__4103\,
            sr => \N__5773\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_43_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5068\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4123\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4629\,
            ce => \N__4103\,
            sr => \N__5773\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_45_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3634\,
            in2 => \_gnd_net_\,
            in3 => \N__5070\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4629\,
            ce => \N__4103\,
            sr => \N__5773\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_17_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5067\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3670\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4629\,
            ce => \N__4103\,
            sr => \N__5773\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_16_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__3676\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5066\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4629\,
            ce => \N__4103\,
            sr => \N__5773\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_6_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__5073\,
            in1 => \N__3664\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4629\,
            ce => \N__4103\,
            sr => \N__5773\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_46_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3652\,
            in2 => \_gnd_net_\,
            in3 => \N__5071\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4629\,
            ce => \N__4103\,
            sr => \N__5773\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_44_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5069\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3640\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4629\,
            ce => \N__4103\,
            sr => \N__5773\
        );

    \fsm_ctrl_inst1.counter_stat_0_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3843\,
            in1 => \N__3742\,
            in2 => \_gnd_net_\,
            in3 => \N__3628\,
            lcout => \fsm_ctrl_inst1.counter_statZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_6_21_0_\,
            carryout => \fsm_ctrl_inst1.counter_stat_cry_0\,
            clk => \N__4625\,
            ce => \N__3799\,
            sr => \N__5775\
        );

    \fsm_ctrl_inst1.counter_stat_1_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3861\,
            in1 => \N__3775\,
            in2 => \_gnd_net_\,
            in3 => \N__3625\,
            lcout => \fsm_ctrl_inst1.counter_statZ0Z_1\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_stat_cry_0\,
            carryout => \fsm_ctrl_inst1.counter_stat_cry_1\,
            clk => \N__4625\,
            ce => \N__3799\,
            sr => \N__5775\
        );

    \fsm_ctrl_inst1.counter_stat_2_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3844\,
            in1 => \N__3711\,
            in2 => \_gnd_net_\,
            in3 => \N__3622\,
            lcout => \fsm_ctrl_inst1.counter_statZ0Z_2\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_stat_cry_1\,
            carryout => \fsm_ctrl_inst1.counter_stat_cry_2\,
            clk => \N__4625\,
            ce => \N__3799\,
            sr => \N__5775\
        );

    \fsm_ctrl_inst1.counter_stat_3_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3862\,
            in1 => \N__3793\,
            in2 => \_gnd_net_\,
            in3 => \N__3874\,
            lcout => \fsm_ctrl_inst1.counter_statZ0Z_3\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_stat_cry_2\,
            carryout => \fsm_ctrl_inst1.counter_stat_cry_3\,
            clk => \N__4625\,
            ce => \N__3799\,
            sr => \N__5775\
        );

    \fsm_ctrl_inst1.counter_stat_4_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3845\,
            in1 => \N__3696\,
            in2 => \_gnd_net_\,
            in3 => \N__3871\,
            lcout => \fsm_ctrl_inst1.counter_statZ0Z_4\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_stat_cry_3\,
            carryout => \fsm_ctrl_inst1.counter_stat_cry_4\,
            clk => \N__4625\,
            ce => \N__3799\,
            sr => \N__5775\
        );

    \fsm_ctrl_inst1.counter_stat_5_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3863\,
            in1 => \N__3729\,
            in2 => \_gnd_net_\,
            in3 => \N__3868\,
            lcout => \fsm_ctrl_inst1.counter_statZ0Z_5\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_stat_cry_4\,
            carryout => \fsm_ctrl_inst1.counter_stat_cry_5\,
            clk => \N__4625\,
            ce => \N__3799\,
            sr => \N__5775\
        );

    \fsm_ctrl_inst1.counter_stat_6_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3846\,
            in1 => \N__3762\,
            in2 => \_gnd_net_\,
            in3 => \N__3802\,
            lcout => \fsm_ctrl_inst1.counter_statZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4625\,
            ce => \N__3799\,
            sr => \N__5775\
        );

    \fsm_ctrl_inst1.current_state_0_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000011101010"
        )
    port map (
            in0 => \N__4760\,
            in1 => \N__4492\,
            in2 => \N__4483\,
            in3 => \N__4311\,
            lcout => \fsm_ctrl_inst1.current_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4624\,
            ce => 'H',
            sr => \N__5778\
        );

    \fsm_ctrl_inst1.current_state_RNO_1_1_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__3791\,
            in1 => \N__3774\,
            in2 => \N__3763\,
            in3 => \N__3741\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.current_state_ns_i_a3_0_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.current_state_RNO_0_1_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__3728\,
            in1 => \N__3712\,
            in2 => \N__3700\,
            in3 => \N__3697\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.current_state_ns_i_a3_0_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.current_state_1_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010111000001100"
        )
    port map (
            in0 => \N__4312\,
            in1 => \N__5033\,
            in2 => \N__3679\,
            in3 => \N__4761\,
            lcout => \fsm_ctrl_inst1.current_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4624\,
            ce => 'H',
            sr => \N__5778\
        );

    \config_register_latched_dec_inst1.DYNSR_0_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4527\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5966\,
            ce => \N__3894\,
            sr => \N__5780\
        );

    \config_register_latched_dec_inst1.DYNSR_1_LC_6_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3943\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5966\,
            ce => \N__3894\,
            sr => \N__5780\
        );

    \config_register_latched_dec_inst1.DYNSR_10_LC_6_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3931\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5966\,
            ce => \N__3894\,
            sr => \N__5780\
        );

    \config_register_latched_dec_inst1.DYNSR_11_LC_6_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3925\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5966\,
            ce => \N__3894\,
            sr => \N__5780\
        );

    \config_register_latched_dec_inst1.DYNSR_12_LC_6_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3919\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5966\,
            ce => \N__3894\,
            sr => \N__5780\
        );

    \config_register_latched_dec_inst1.DYNSR_13_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3913\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5966\,
            ce => \N__3894\,
            sr => \N__5780\
        );

    \config_register_latched_dec_inst1.DYNSR_14_LC_6_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3907\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5966\,
            ce => \N__3894\,
            sr => \N__5780\
        );

    \config_register_latched_dec_inst1.DYNSR_15_LC_6_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3901\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5966\,
            ce => \N__3894\,
            sr => \N__5780\
        );

    \config_register_latched_dec_inst1.DYNSR_cnv_0_LC_6_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__4230\,
            in1 => \N__4022\,
            in2 => \_gnd_net_\,
            in3 => \N__4006\,
            lcout => \config_register_latched_dec_inst1.DYNSR_cnvZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.CLK_uC_0_LC_6_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4023\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_ctrl_inst1_CLK_uC_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5967\,
            ce => 'H',
            sr => \N__5782\
        );

    \fsm_ctrl_inst1.toggle_clk_uC4_0_LC_6_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4339\,
            lcout => \toggle_clk_uC4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5968\,
            ce => 'H',
            sr => \N__5784\
        );

    \config_register_latched_dec_inst1.STATSR_cnv_0_LC_6_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__4234\,
            in1 => \_gnd_net_\,
            in2 => \N__4024\,
            in3 => \N__4005\,
            lcout => \STATSR_cnv_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_RNIMLJF1_4_LC_6_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4409\,
            in1 => \N__4451\,
            in2 => \N__4366\,
            in3 => \N__4430\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.counter_idlelde_0_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.current_state_RNIPMA12_0_LC_6_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5048\,
            in2 => \N__3976\,
            in3 => \N__4772\,
            lcout => \fsm_ctrl_inst1.counter_idlee_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_79_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3973\,
            in2 => \_gnd_net_\,
            in3 => \N__5168\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4635\,
            ce => \N__4102\,
            sr => \N__5770\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_52_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4162\,
            in2 => \_gnd_net_\,
            in3 => \N__5116\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4630\,
            ce => \N__4104\,
            sr => \N__5774\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_38_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5113\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4174\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4630\,
            ce => \N__4104\,
            sr => \N__5774\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_36_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3955\,
            in2 => \_gnd_net_\,
            in3 => \N__5111\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4630\,
            ce => \N__4104\,
            sr => \N__5774\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_50_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5114\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3949\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4630\,
            ce => \N__4104\,
            sr => \N__5774\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_37_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4180\,
            in2 => \_gnd_net_\,
            in3 => \N__5112\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4630\,
            ce => \N__4104\,
            sr => \N__5774\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_51_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5115\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4168\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4630\,
            ce => \N__4104\,
            sr => \N__5774\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_40_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5107\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4150\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4626\,
            ce => \N__4105\,
            sr => \N__5776\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_39_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4156\,
            in2 => \_gnd_net_\,
            in3 => \N__5106\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4626\,
            ce => \N__4105\,
            sr => \N__5776\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_87_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5110\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4144\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4626\,
            ce => \N__4105\,
            sr => \N__5776\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_18_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4138\,
            in2 => \_gnd_net_\,
            in3 => \N__5105\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4626\,
            ce => \N__4105\,
            sr => \N__5776\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_42_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5109\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4111\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4626\,
            ce => \N__4105\,
            sr => \N__5776\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_41_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4117\,
            in2 => \_gnd_net_\,
            in3 => \N__5108\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4626\,
            ce => \N__4105\,
            sr => \N__5776\
        );

    \fsm_ctrl_inst1.current_state_RNI1GR8_0_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4729\,
            lcout => \fsm_ctrl_inst1.current_state_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.SEL_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4767\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \SEL_REG\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4622\,
            ce => 'H',
            sr => \N__5781\
        );

    \fsm_ctrl_inst1.MOSI_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__4333\,
            in1 => \N__4766\,
            in2 => \N__4324\,
            in3 => \N__5034\,
            lcout => \MOSI\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4622\,
            ce => 'H',
            sr => \N__5781\
        );

    \fsm_ctrl_inst1.counter_din_RNI6L3H1_3_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4280\,
            in1 => \N__4246\,
            in2 => \N__4299\,
            in3 => \N__4266\,
            lcout => \fsm_ctrl_inst1.N_119_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_din_0_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__4268\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4763\,
            lcout => \fsm_ctrl_inst1.counter_dinZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4621\,
            ce => 'H',
            sr => \N__5783\
        );

    \fsm_ctrl_inst1.counter_din_RNO_0_3_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__4281\,
            in1 => \N__4247\,
            in2 => \N__4300\,
            in3 => \N__4267\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.N_105_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_din_3_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4303\,
            in3 => \N__4764\,
            lcout => \fsm_ctrl_inst1.counter_dinZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4621\,
            ce => 'H',
            sr => \N__5783\
        );

    \fsm_ctrl_inst1.counter_din_2_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010100010100000"
        )
    port map (
            in0 => \N__4762\,
            in1 => \N__4251\,
            in2 => \N__4285\,
            in3 => \N__4270\,
            lcout => \fsm_ctrl_inst1.counter_dinZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4621\,
            ce => 'H',
            sr => \N__5783\
        );

    \fsm_ctrl_inst1.counter_din_1_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__4269\,
            in1 => \_gnd_net_\,
            in2 => \N__4252\,
            in3 => \N__4765\,
            lcout => \fsm_ctrl_inst1.counter_dinZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4621\,
            ce => 'H',
            sr => \N__5783\
        );

    \config_register_latched_dec_inst1.DYNSR_RNIQ2U9_15_LC_7_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4223\,
            in1 => \N__4210\,
            in2 => \_gnd_net_\,
            in3 => \N__4543\,
            lcout => \SDO_signal_out_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.current_state_RNO_1_0_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__5036\,
            in1 => \N__4453\,
            in2 => \N__4471\,
            in3 => \N__4364\,
            lcout => \fsm_ctrl_inst1.current_state_ns_0_i_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.current_state_RNO_0_0_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4410\,
            in2 => \_gnd_net_\,
            in3 => \N__4431\,
            lcout => \fsm_ctrl_inst1.N_122_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.current_state_RNI31NH_0_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__5035\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4768\,
            lcout => \fsm_ctrl_inst1.current_state_23_d_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_0_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4389\,
            in1 => \N__4467\,
            in2 => \_gnd_net_\,
            in3 => \N__4456\,
            lcout => \fsm_ctrl_inst1.counter_idleZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_25_0_\,
            carryout => \fsm_ctrl_inst1.counter_idle_cry_0\,
            clk => \N__4620\,
            ce => \N__4345\,
            sr => \N__5785\
        );

    \fsm_ctrl_inst1.counter_idle_1_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4386\,
            in1 => \N__4452\,
            in2 => \_gnd_net_\,
            in3 => \N__4435\,
            lcout => \fsm_ctrl_inst1.counter_idleZ0Z_1\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_idle_cry_0\,
            carryout => \fsm_ctrl_inst1.counter_idle_cry_1\,
            clk => \N__4620\,
            ce => \N__4345\,
            sr => \N__5785\
        );

    \fsm_ctrl_inst1.counter_idle_2_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4390\,
            in1 => \N__4432\,
            in2 => \_gnd_net_\,
            in3 => \N__4414\,
            lcout => \fsm_ctrl_inst1.counter_idleZ0Z_2\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_idle_cry_1\,
            carryout => \fsm_ctrl_inst1.counter_idle_cry_2\,
            clk => \N__4620\,
            ce => \N__4345\,
            sr => \N__5785\
        );

    \fsm_ctrl_inst1.counter_idle_3_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4387\,
            in1 => \N__4411\,
            in2 => \_gnd_net_\,
            in3 => \N__4393\,
            lcout => \fsm_ctrl_inst1.counter_idleZ0Z_3\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_idle_cry_2\,
            carryout => \fsm_ctrl_inst1.counter_idle_cry_3\,
            clk => \N__4620\,
            ce => \N__4345\,
            sr => \N__5785\
        );

    \fsm_ctrl_inst1.counter_idle_4_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__4365\,
            in1 => \N__4388\,
            in2 => \_gnd_net_\,
            in3 => \N__4369\,
            lcout => \fsm_ctrl_inst1.counter_idleZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4620\,
            ce => \N__4345\,
            sr => \N__5785\
        );

    \fsm_ctrl_inst1.toggle_clk_uC3_0_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5197\,
            lcout => \fsm_ctrl_inst1.toggle_clk_uC3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5970\,
            ce => 'H',
            sr => \N__5787\
        );

    \fsm_ctrl_inst1.toggle_clk_uC2_0_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4552\,
            lcout => \fsm_ctrl_inst1.toggle_clk_uC2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5970\,
            ce => 'H',
            sr => \N__5787\
        );

    \fsm_ctrl_inst1.toggle_clk_uC1_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__5191\,
            in1 => \N__4551\,
            in2 => \N__4780\,
            in3 => \N__4651\,
            lcout => \fsm_ctrl_inst1.toggle_clk_uCZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5970\,
            ce => 'H',
            sr => \N__5787\
        );

    \config_register_latched_dec_inst1.STATSR_87_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4510\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5969\,
            ce => \N__5896\,
            sr => \N__5786\
        );

    \config_register_latched_dec_inst1.STATSR_0_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4534\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5971\,
            ce => \N__5895\,
            sr => \N__5788\
        );

    \config_register_latched_dec_inst1.STATSR_85_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5239\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5971\,
            ce => \N__5895\,
            sr => \N__5788\
        );

    \config_register_latched_dec_inst1.STATSR_86_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4516\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5971\,
            ce => \N__5895\,
            sr => \N__5788\
        );

    \config_register_latched_dec_inst1.STATSR_3_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5245\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5972\,
            ce => \N__5894\,
            sr => \N__5789\
        );

    \config_register_latched_dec_inst1.STATSR_1_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4504\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5972\,
            ce => \N__5894\,
            sr => \N__5789\
        );

    \config_register_latched_dec_inst1.STATSR_4_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4498\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5972\,
            ce => \N__5894\,
            sr => \N__5789\
        );

    \config_register_latched_dec_inst1.STATSR_2_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5251\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5972\,
            ce => \N__5894\,
            sr => \N__5789\
        );

    \config_register_latched_dec_inst1.STATSR_84_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5233\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5972\,
            ce => \N__5894\,
            sr => \N__5789\
        );

    \config_register_latched_dec_inst1.STATSR_83_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5215\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5973\,
            ce => \N__5893\,
            sr => \N__5790\
        );

    \config_register_latched_dec_inst1.STATSR_5_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5227\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5973\,
            ce => \N__5893\,
            sr => \N__5790\
        );

    \config_register_latched_dec_inst1.STATSR_6_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5221\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5974\,
            ce => \N__5892\,
            sr => \N__5791\
        );

    \config_register_latched_dec_inst1.STATSR_82_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5269\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5974\,
            ce => \N__5892\,
            sr => \N__5791\
        );

    \config_register_latched_dec_inst1.STATSR_7_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5209\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5975\,
            ce => \N__5890\,
            sr => \N__5792\
        );

    \config_register_latched_dec_inst1.STATSR_8_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5203\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5977\,
            ce => \N__5888\,
            sr => \N__5794\
        );

    \config_register_latched_dec_inst1.STATSR_10_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5299\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5979\,
            ce => \N__5887\,
            sr => \N__5796\
        );

    \config_register_latched_dec_inst1.STATSR_9_LC_12_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5305\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5979\,
            ce => \N__5887\,
            sr => \N__5796\
        );

    \config_register_latched_dec_inst1.STATSR_12_LC_12_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5287\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5979\,
            ce => \N__5887\,
            sr => \N__5796\
        );

    \config_register_latched_dec_inst1.STATSR_11_LC_12_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5293\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5979\,
            ce => \N__5887\,
            sr => \N__5796\
        );

    \config_register_latched_dec_inst1.STATSR_79_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5263\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5976\,
            ce => \N__5891\,
            sr => \N__5793\
        );

    \config_register_latched_dec_inst1.STATSR_80_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5281\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5976\,
            ce => \N__5891\,
            sr => \N__5793\
        );

    \config_register_latched_dec_inst1.STATSR_81_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5275\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5976\,
            ce => \N__5891\,
            sr => \N__5793\
        );

    \config_register_latched_dec_inst1.STATSR_78_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5257\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5978\,
            ce => \N__5889\,
            sr => \N__5795\
        );

    \config_register_latched_dec_inst1.STATSR_77_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5323\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5978\,
            ce => \N__5889\,
            sr => \N__5795\
        );

    \config_register_latched_dec_inst1.STATSR_15_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5359\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5980\,
            ce => \N__5885\,
            sr => \N__5797\
        );

    \config_register_latched_dec_inst1.STATSR_14_LC_13_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5347\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5980\,
            ce => \N__5885\,
            sr => \N__5797\
        );

    \config_register_latched_dec_inst1.STATSR_13_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5353\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5980\,
            ce => \N__5885\,
            sr => \N__5797\
        );

    \config_register_latched_dec_inst1.STATSR_16_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5341\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5980\,
            ce => \N__5885\,
            sr => \N__5797\
        );

    \config_register_latched_dec_inst1.STATSR_74_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5317\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5981\,
            ce => \N__5886\,
            sr => \N__5798\
        );

    \config_register_latched_dec_inst1.STATSR_75_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5335\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5981\,
            ce => \N__5886\,
            sr => \N__5798\
        );

    \config_register_latched_dec_inst1.STATSR_76_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5329\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5981\,
            ce => \N__5886\,
            sr => \N__5798\
        );

    \config_register_latched_dec_inst1.STATSR_73_LC_14_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5407\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5982\,
            ce => \N__5884\,
            sr => \N__5799\
        );

    \config_register_latched_dec_inst1.STATSR_17_LC_14_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5311\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5982\,
            ce => \N__5884\,
            sr => \N__5799\
        );

    \config_register_latched_dec_inst1.STATSR_69_LC_14_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5401\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5983\,
            ce => \N__5882\,
            sr => \N__5800\
        );

    \config_register_latched_dec_inst1.STATSR_71_LC_14_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5389\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5983\,
            ce => \N__5882\,
            sr => \N__5800\
        );

    \config_register_latched_dec_inst1.STATSR_72_LC_14_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5413\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5983\,
            ce => \N__5882\,
            sr => \N__5800\
        );

    \config_register_latched_dec_inst1.STATSR_68_LC_14_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5377\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5983\,
            ce => \N__5882\,
            sr => \N__5800\
        );

    \config_register_latched_dec_inst1.STATSR_70_LC_14_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5395\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5983\,
            ce => \N__5882\,
            sr => \N__5800\
        );

    \config_register_latched_dec_inst1.STATSR_66_LC_14_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5371\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5983\,
            ce => \N__5882\,
            sr => \N__5800\
        );

    \config_register_latched_dec_inst1.STATSR_67_LC_14_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5383\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5983\,
            ce => \N__5882\,
            sr => \N__5800\
        );

    \config_register_latched_dec_inst1.STATSR_65_LC_14_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5461\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5985\,
            ce => \N__5879\,
            sr => \N__5802\
        );

    \config_register_latched_dec_inst1.STATSR_63_LC_14_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5365\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5985\,
            ce => \N__5879\,
            sr => \N__5802\
        );

    \config_register_latched_dec_inst1.STATSR_62_LC_14_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5473\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5985\,
            ce => \N__5879\,
            sr => \N__5802\
        );

    \config_register_latched_dec_inst1.STATSR_61_LC_14_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5437\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5985\,
            ce => \N__5879\,
            sr => \N__5802\
        );

    \config_register_latched_dec_inst1.STATSR_64_LC_14_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5467\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5985\,
            ce => \N__5879\,
            sr => \N__5802\
        );

    \config_register_latched_dec_inst1.STATSR_18_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5455\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5984\,
            ce => \N__5883\,
            sr => \N__5801\
        );

    \config_register_latched_dec_inst1.STATSR_19_LC_15_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5449\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5984\,
            ce => \N__5883\,
            sr => \N__5801\
        );

    \config_register_latched_dec_inst1.STATSR_56_LC_15_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5503\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5986\,
            ce => \N__5880\,
            sr => \N__5803\
        );

    \config_register_latched_dec_inst1.STATSR_57_LC_15_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5443\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5988\,
            ce => \N__5877\,
            sr => \N__5805\
        );

    \config_register_latched_dec_inst1.STATSR_60_LC_15_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5419\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5988\,
            ce => \N__5877\,
            sr => \N__5805\
        );

    \config_register_latched_dec_inst1.STATSR_58_LC_15_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5431\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5988\,
            ce => \N__5877\,
            sr => \N__5805\
        );

    \config_register_latched_dec_inst1.STATSR_59_LC_15_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5425\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5988\,
            ce => \N__5877\,
            sr => \N__5805\
        );

    \config_register_latched_dec_inst1.STATSR_51_LC_16_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5527\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5987\,
            ce => \N__5881\,
            sr => \N__5804\
        );

    \config_register_latched_dec_inst1.STATSR_50_LC_16_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5521\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5987\,
            ce => \N__5881\,
            sr => \N__5804\
        );

    \config_register_latched_dec_inst1.STATSR_49_LC_16_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5599\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5987\,
            ce => \N__5881\,
            sr => \N__5804\
        );

    \config_register_latched_dec_inst1.STATSR_54_LC_16_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5515\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5989\,
            ce => \N__5878\,
            sr => \N__5806\
        );

    \config_register_latched_dec_inst1.STATSR_53_LC_16_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5491\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5989\,
            ce => \N__5878\,
            sr => \N__5806\
        );

    \config_register_latched_dec_inst1.STATSR_55_LC_16_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5509\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5989\,
            ce => \N__5878\,
            sr => \N__5806\
        );

    \config_register_latched_dec_inst1.STATSR_52_LC_16_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5497\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5989\,
            ce => \N__5878\,
            sr => \N__5806\
        );

    \config_register_latched_dec_inst1.STATSR_20_LC_16_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5485\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5989\,
            ce => \N__5878\,
            sr => \N__5806\
        );

    \config_register_latched_dec_inst1.STATSR_21_LC_16_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5479\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5991\,
            ce => \N__5875\,
            sr => \N__5808\
        );

    \config_register_latched_dec_inst1.STATSR_35_LC_16_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5575\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5991\,
            ce => \N__5875\,
            sr => \N__5808\
        );

    \config_register_latched_dec_inst1.STATSR_33_LC_16_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5539\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5991\,
            ce => \N__5875\,
            sr => \N__5808\
        );

    \config_register_latched_dec_inst1.STATSR_34_LC_16_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5581\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5991\,
            ce => \N__5875\,
            sr => \N__5808\
        );

    \config_register_latched_dec_inst1.STATSR_22_LC_16_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5569\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5993\,
            ce => \N__5873\,
            sr => \N__5810\
        );

    \config_register_latched_dec_inst1.STATSR_24_LC_16_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5551\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5993\,
            ce => \N__5873\,
            sr => \N__5810\
        );

    \config_register_latched_dec_inst1.STATSR_30_LC_16_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5617\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5993\,
            ce => \N__5873\,
            sr => \N__5810\
        );

    \config_register_latched_dec_inst1.STATSR_31_LC_16_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5563\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5993\,
            ce => \N__5873\,
            sr => \N__5810\
        );

    \config_register_latched_dec_inst1.STATSR_23_LC_16_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5557\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5993\,
            ce => \N__5873\,
            sr => \N__5810\
        );

    \config_register_latched_dec_inst1.STATSR_32_LC_16_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5545\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5993\,
            ce => \N__5873\,
            sr => \N__5810\
        );

    \config_register_latched_dec_inst1.STATSR_25_LC_16_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5533\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5995\,
            ce => \N__5871\,
            sr => \N__5812\
        );

    \config_register_latched_dec_inst1.STATSR_27_LC_16_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5623\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5995\,
            ce => \N__5871\,
            sr => \N__5812\
        );

    \config_register_latched_dec_inst1.STATSR_26_LC_16_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5629\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5995\,
            ce => \N__5871\,
            sr => \N__5812\
        );

    \config_register_latched_dec_inst1.STATSR_29_LC_16_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5605\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5995\,
            ce => \N__5871\,
            sr => \N__5812\
        );

    \config_register_latched_dec_inst1.STATSR_28_LC_16_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5611\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5995\,
            ce => \N__5871\,
            sr => \N__5812\
        );

    \config_register_latched_dec_inst1.STATSR_48_LC_17_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6043\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5990\,
            ce => \N__5876\,
            sr => \N__5807\
        );

    \config_register_latched_dec_inst1.STATSR_43_LC_17_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5593\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5990\,
            ce => \N__5876\,
            sr => \N__5807\
        );

    \config_register_latched_dec_inst1.STATSR_46_LC_17_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6055\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5990\,
            ce => \N__5876\,
            sr => \N__5807\
        );

    \config_register_latched_dec_inst1.STATSR_42_LC_17_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6037\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5990\,
            ce => \N__5876\,
            sr => \N__5807\
        );

    \config_register_latched_dec_inst1.STATSR_44_LC_17_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5587\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5990\,
            ce => \N__5876\,
            sr => \N__5807\
        );

    \config_register_latched_dec_inst1.STATSR_45_LC_17_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6061\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5990\,
            ce => \N__5876\,
            sr => \N__5807\
        );

    \config_register_latched_dec_inst1.STATSR_47_LC_17_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6049\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5990\,
            ce => \N__5876\,
            sr => \N__5807\
        );

    \config_register_latched_dec_inst1.STATSR_41_LC_17_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6031\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5992\,
            ce => \N__5874\,
            sr => \N__5809\
        );

    \config_register_latched_dec_inst1.STATSR_40_LC_17_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6019\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5992\,
            ce => \N__5874\,
            sr => \N__5809\
        );

    \config_register_latched_dec_inst1.STATSR_38_LC_17_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6001\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5992\,
            ce => \N__5874\,
            sr => \N__5809\
        );

    \config_register_latched_dec_inst1.STATSR_39_LC_17_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6025\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5992\,
            ce => \N__5874\,
            sr => \N__5809\
        );

    \config_register_latched_dec_inst1.STATSR_36_LC_17_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6013\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5994\,
            ce => \N__5872\,
            sr => \N__5811\
        );

    \config_register_latched_dec_inst1.STATSR_37_LC_17_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6007\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5994\,
            ce => \N__5872\,
            sr => \N__5811\
        );
end \INTERFACE\;
