// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 13 2025 09:52:51

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    signal_out,
    CLK,
    SELSTAT,
    SELDYN,
    RST_N);

    output signal_out;
    input CLK;
    input SELSTAT;
    input SELDYN;
    input RST_N;

    wire N__2717;
    wire N__2716;
    wire N__2715;
    wire N__2706;
    wire N__2705;
    wire N__2704;
    wire N__2697;
    wire N__2696;
    wire N__2695;
    wire N__2688;
    wire N__2687;
    wire N__2686;
    wire N__2679;
    wire N__2678;
    wire N__2677;
    wire N__2660;
    wire N__2657;
    wire N__2654;
    wire N__2651;
    wire N__2648;
    wire N__2645;
    wire N__2642;
    wire N__2639;
    wire N__2636;
    wire N__2633;
    wire N__2630;
    wire N__2627;
    wire N__2624;
    wire N__2621;
    wire N__2618;
    wire N__2615;
    wire N__2612;
    wire N__2611;
    wire N__2610;
    wire N__2609;
    wire N__2608;
    wire N__2607;
    wire N__2606;
    wire N__2605;
    wire N__2604;
    wire N__2603;
    wire N__2602;
    wire N__2601;
    wire N__2600;
    wire N__2599;
    wire N__2598;
    wire N__2597;
    wire N__2596;
    wire N__2595;
    wire N__2594;
    wire N__2593;
    wire N__2592;
    wire N__2591;
    wire N__2590;
    wire N__2589;
    wire N__2588;
    wire N__2587;
    wire N__2586;
    wire N__2585;
    wire N__2584;
    wire N__2583;
    wire N__2582;
    wire N__2581;
    wire N__2580;
    wire N__2579;
    wire N__2578;
    wire N__2577;
    wire N__2576;
    wire N__2575;
    wire N__2574;
    wire N__2573;
    wire N__2572;
    wire N__2571;
    wire N__2570;
    wire N__2569;
    wire N__2568;
    wire N__2567;
    wire N__2566;
    wire N__2565;
    wire N__2560;
    wire N__2549;
    wire N__2540;
    wire N__2539;
    wire N__2538;
    wire N__2537;
    wire N__2536;
    wire N__2535;
    wire N__2534;
    wire N__2533;
    wire N__2532;
    wire N__2531;
    wire N__2530;
    wire N__2529;
    wire N__2528;
    wire N__2527;
    wire N__2526;
    wire N__2515;
    wire N__2500;
    wire N__2491;
    wire N__2476;
    wire N__2459;
    wire N__2446;
    wire N__2443;
    wire N__2438;
    wire N__2425;
    wire N__2408;
    wire N__2395;
    wire N__2386;
    wire N__2385;
    wire N__2384;
    wire N__2383;
    wire N__2382;
    wire N__2381;
    wire N__2380;
    wire N__2379;
    wire N__2378;
    wire N__2377;
    wire N__2376;
    wire N__2375;
    wire N__2374;
    wire N__2373;
    wire N__2372;
    wire N__2371;
    wire N__2370;
    wire N__2369;
    wire N__2368;
    wire N__2367;
    wire N__2366;
    wire N__2365;
    wire N__2364;
    wire N__2361;
    wire N__2358;
    wire N__2345;
    wire N__2328;
    wire N__2327;
    wire N__2326;
    wire N__2325;
    wire N__2324;
    wire N__2323;
    wire N__2322;
    wire N__2305;
    wire N__2296;
    wire N__2283;
    wire N__2276;
    wire N__2273;
    wire N__2270;
    wire N__2267;
    wire N__2264;
    wire N__2263;
    wire N__2262;
    wire N__2261;
    wire N__2260;
    wire N__2259;
    wire N__2258;
    wire N__2257;
    wire N__2256;
    wire N__2255;
    wire N__2254;
    wire N__2253;
    wire N__2252;
    wire N__2251;
    wire N__2250;
    wire N__2249;
    wire N__2248;
    wire N__2213;
    wire N__2210;
    wire N__2207;
    wire N__2206;
    wire N__2205;
    wire N__2204;
    wire N__2203;
    wire N__2202;
    wire N__2201;
    wire N__2200;
    wire N__2199;
    wire N__2198;
    wire N__2197;
    wire N__2196;
    wire N__2195;
    wire N__2194;
    wire N__2165;
    wire N__2162;
    wire N__2159;
    wire N__2158;
    wire N__2157;
    wire N__2156;
    wire N__2155;
    wire N__2154;
    wire N__2153;
    wire N__2152;
    wire N__2151;
    wire N__2150;
    wire N__2149;
    wire N__2148;
    wire N__2147;
    wire N__2146;
    wire N__2145;
    wire N__2144;
    wire N__2143;
    wire N__2108;
    wire N__2105;
    wire N__2102;
    wire N__2099;
    wire N__2096;
    wire N__2093;
    wire N__2090;
    wire N__2087;
    wire N__2084;
    wire N__2081;
    wire N__2078;
    wire N__2075;
    wire N__2072;
    wire N__2069;
    wire N__2066;
    wire N__2063;
    wire N__2060;
    wire N__2057;
    wire N__2054;
    wire N__2051;
    wire N__2048;
    wire N__2045;
    wire N__2042;
    wire N__2039;
    wire N__2036;
    wire N__2033;
    wire N__2030;
    wire N__2027;
    wire N__2024;
    wire N__2021;
    wire N__2018;
    wire N__2015;
    wire N__2012;
    wire N__2009;
    wire N__2006;
    wire N__2003;
    wire N__2000;
    wire N__1997;
    wire N__1994;
    wire N__1991;
    wire N__1988;
    wire N__1985;
    wire N__1982;
    wire N__1979;
    wire N__1976;
    wire N__1973;
    wire N__1970;
    wire N__1967;
    wire N__1964;
    wire N__1961;
    wire N__1958;
    wire N__1955;
    wire N__1952;
    wire N__1949;
    wire N__1946;
    wire N__1943;
    wire N__1940;
    wire N__1937;
    wire N__1934;
    wire N__1931;
    wire N__1928;
    wire N__1925;
    wire N__1922;
    wire N__1919;
    wire N__1916;
    wire N__1913;
    wire N__1910;
    wire N__1907;
    wire N__1904;
    wire N__1901;
    wire N__1898;
    wire N__1895;
    wire N__1892;
    wire N__1889;
    wire N__1886;
    wire N__1883;
    wire N__1880;
    wire N__1877;
    wire N__1874;
    wire N__1871;
    wire N__1868;
    wire N__1865;
    wire N__1862;
    wire N__1859;
    wire N__1856;
    wire N__1853;
    wire N__1850;
    wire N__1847;
    wire N__1844;
    wire N__1841;
    wire N__1838;
    wire N__1835;
    wire N__1832;
    wire N__1829;
    wire N__1826;
    wire N__1823;
    wire N__1820;
    wire N__1817;
    wire N__1814;
    wire N__1811;
    wire N__1808;
    wire N__1805;
    wire N__1802;
    wire N__1799;
    wire N__1796;
    wire N__1793;
    wire N__1790;
    wire N__1789;
    wire N__1788;
    wire N__1787;
    wire N__1786;
    wire N__1785;
    wire N__1784;
    wire N__1783;
    wire N__1782;
    wire N__1781;
    wire N__1780;
    wire N__1779;
    wire N__1778;
    wire N__1777;
    wire N__1776;
    wire N__1775;
    wire N__1774;
    wire N__1773;
    wire N__1772;
    wire N__1769;
    wire N__1764;
    wire N__1747;
    wire N__1730;
    wire N__1721;
    wire N__1718;
    wire N__1715;
    wire N__1712;
    wire N__1709;
    wire N__1706;
    wire N__1703;
    wire N__1700;
    wire N__1697;
    wire N__1694;
    wire N__1691;
    wire N__1688;
    wire N__1685;
    wire N__1682;
    wire N__1679;
    wire N__1676;
    wire N__1673;
    wire N__1670;
    wire N__1667;
    wire N__1664;
    wire N__1661;
    wire N__1658;
    wire N__1655;
    wire N__1652;
    wire N__1649;
    wire N__1646;
    wire N__1643;
    wire N__1640;
    wire N__1637;
    wire N__1634;
    wire N__1631;
    wire N__1628;
    wire N__1625;
    wire N__1622;
    wire N__1619;
    wire N__1616;
    wire N__1613;
    wire N__1610;
    wire N__1607;
    wire N__1604;
    wire N__1601;
    wire N__1598;
    wire N__1595;
    wire N__1592;
    wire N__1589;
    wire N__1586;
    wire N__1583;
    wire N__1580;
    wire N__1577;
    wire N__1574;
    wire N__1571;
    wire N__1568;
    wire N__1565;
    wire N__1562;
    wire N__1559;
    wire N__1556;
    wire N__1553;
    wire N__1550;
    wire N__1547;
    wire N__1544;
    wire N__1541;
    wire N__1538;
    wire N__1535;
    wire N__1532;
    wire N__1529;
    wire N__1526;
    wire N__1523;
    wire N__1520;
    wire N__1517;
    wire N__1514;
    wire N__1511;
    wire N__1508;
    wire N__1505;
    wire N__1502;
    wire N__1499;
    wire N__1496;
    wire N__1493;
    wire N__1490;
    wire N__1487;
    wire N__1484;
    wire N__1481;
    wire N__1478;
    wire N__1475;
    wire N__1472;
    wire N__1469;
    wire N__1466;
    wire N__1463;
    wire N__1460;
    wire N__1457;
    wire N__1454;
    wire N__1451;
    wire N__1448;
    wire N__1445;
    wire N__1442;
    wire N__1439;
    wire N__1438;
    wire N__1435;
    wire N__1432;
    wire N__1427;
    wire N__1424;
    wire N__1421;
    wire N__1418;
    wire N__1415;
    wire N__1412;
    wire N__1409;
    wire N__1406;
    wire N__1403;
    wire N__1400;
    wire N__1397;
    wire N__1394;
    wire N__1391;
    wire N__1388;
    wire N__1385;
    wire N__1382;
    wire GNDG0;
    wire VCCG0;
    wire \generator_inst1.REGDYNZ0Z_1 ;
    wire \generator_inst1.REGDYNZ0Z_2 ;
    wire \generator_inst1.REGDYNZ0Z_5 ;
    wire \generator_inst1.REGDYNZ0Z_6 ;
    wire \generator_inst1.REGDYNZ0Z_3 ;
    wire \generator_inst1.REGDYNZ0Z_4 ;
    wire \generator_inst1.REGDYNZ0Z_0 ;
    wire \generator_inst1.REGDYNZ0Z_10 ;
    wire \generator_inst1.REGDYNZ0Z_11 ;
    wire \generator_inst1.REGDYNZ0Z_12 ;
    wire \generator_inst1.REGDYNZ0Z_13 ;
    wire \generator_inst1.REGDYNZ0Z_14 ;
    wire \generator_inst1.REGDYNZ0Z_9 ;
    wire \generator_inst1.REGDYNZ0Z_7 ;
    wire \generator_inst1.REGDYNZ0Z_8 ;
    wire \generator_inst1.REGDYNZ0Z_15 ;
    wire generated_signal;
    wire signal_out_c;
    wire \generator_inst1.REGDYN8_iZ0 ;
    wire \generator_inst1.REGSTATZ0Z_86 ;
    wire \generator_inst1.REGSTATZ0Z_87 ;
    wire \generator_inst1.REGSTATZ0Z_84 ;
    wire \generator_inst1.REGSTATZ0Z_85 ;
    wire \generator_inst1.REGSTATZ0Z_9 ;
    wire \generator_inst1.REGSTATZ0Z_6 ;
    wire \generator_inst1.REGSTATZ0Z_7 ;
    wire \generator_inst1.REGSTATZ0Z_8 ;
    wire \generator_inst1.REGSTATZ0Z_10 ;
    wire \generator_inst1.REGSTATZ0Z_11 ;
    wire \generator_inst1.REGSTATZ0Z_12 ;
    wire \generator_inst1.REGSTATZ0Z_13 ;
    wire \generator_inst1.REGSTATZ0Z_18 ;
    wire \generator_inst1.REGSTATZ0Z_14 ;
    wire \generator_inst1.REGSTATZ0Z_15 ;
    wire \generator_inst1.REGSTATZ0Z_16 ;
    wire \generator_inst1.REGSTATZ0Z_17 ;
    wire \generator_inst1.REGSTATZ0Z_34 ;
    wire \generator_inst1.REGSTATZ0Z_35 ;
    wire \generator_inst1.REGSTATZ0Z_36 ;
    wire \generator_inst1.REGSTATZ0Z_32 ;
    wire \generator_inst1.REGSTATZ0Z_33 ;
    wire \generator_inst1.REGSTATZ0Z_37 ;
    wire \generator_inst1.REGSTATZ0Z_38 ;
    wire \generator_inst1.REGSTATZ0Z_39 ;
    wire \generator_inst1.REGSTATZ0Z_40 ;
    wire \generator_inst1.REGSTATZ0Z_41 ;
    wire \generator_inst1.REGSTATZ0Z_42 ;
    wire \generator_inst1.REGSTATZ0Z_43 ;
    wire \generator_inst1.REGSTATZ0Z_44 ;
    wire SELDYN_c;
    wire SELDYN_c_i;
    wire RST_N_c;
    wire RST_N_c_i;
    wire \generator_inst1.REGSTATZ0Z_80 ;
    wire \generator_inst1.REGSTATZ0Z_81 ;
    wire \generator_inst1.REGSTATZ0Z_79 ;
    wire \generator_inst1.REGSTATZ0Z_82 ;
    wire \generator_inst1.REGSTATZ0Z_83 ;
    wire \generator_inst1.REGSTATZ0Z_5 ;
    wire \generator_inst1.REGSTATZ0Z_2 ;
    wire \generator_inst1.REGSTATZ0Z_3 ;
    wire \generator_inst1.REGSTATZ0Z_4 ;
    wire \generator_inst1.REGSTATZ0Z_24 ;
    wire \generator_inst1.REGSTATZ0Z_23 ;
    wire \generator_inst1.REGSTATZ0Z_19 ;
    wire \generator_inst1.REGSTATZ0Z_22 ;
    wire \generator_inst1.REGSTATZ0Z_20 ;
    wire \generator_inst1.REGSTATZ0Z_21 ;
    wire \generator_inst1.REGSTATZ0Z_0 ;
    wire \generator_inst1.REGSTATZ0Z_1 ;
    wire \generator_inst1.REGSTATZ0Z_27 ;
    wire \generator_inst1.REGSTATZ0Z_28 ;
    wire \generator_inst1.REGSTATZ0Z_29 ;
    wire \generator_inst1.REGSTATZ0Z_25 ;
    wire \generator_inst1.REGSTATZ0Z_26 ;
    wire \generator_inst1.REGSTATZ0Z_30 ;
    wire \generator_inst1.REGSTATZ0Z_31 ;
    wire \generator_inst1.REGSTATZ0Z_51 ;
    wire \generator_inst1.REGSTATZ0Z_52 ;
    wire \generator_inst1.REGSTATZ0Z_45 ;
    wire \generator_inst1.REGSTATZ0Z_46 ;
    wire \generator_inst1.REGSTATZ0Z_47 ;
    wire \generator_inst1.REGSTATZ0Z_48 ;
    wire \generator_inst1.REGSTATZ0Z_49 ;
    wire \generator_inst1.REGSTATZ0Z_50 ;
    wire \generator_inst1.REGSTATZ0Z_76 ;
    wire \generator_inst1.REGSTATZ0Z_77 ;
    wire \generator_inst1.REGSTATZ0Z_78 ;
    wire \generator_inst1.REGSTATZ0Z_75 ;
    wire \generator_inst1.REGSTATZ0Z_74 ;
    wire \generator_inst1.REGSTATZ0Z_73 ;
    wire \generator_inst1.REGSTATZ0Z_67 ;
    wire \generator_inst1.REGSTATZ0Z_70 ;
    wire \generator_inst1.REGSTATZ0Z_68 ;
    wire \generator_inst1.REGSTATZ0Z_69 ;
    wire \generator_inst1.REGSTATZ0Z_71 ;
    wire \generator_inst1.REGSTATZ0Z_72 ;
    wire \generator_inst1.REGSTATZ0Z_63 ;
    wire \generator_inst1.REGSTATZ0Z_62 ;
    wire \generator_inst1.REGSTATZ0Z_60 ;
    wire \generator_inst1.REGSTATZ0Z_61 ;
    wire \generator_inst1.REGSTATZ0Z_66 ;
    wire \generator_inst1.REGSTATZ0Z_64 ;
    wire \generator_inst1.REGSTATZ0Z_65 ;
    wire \generator_inst1.REGSTATZ0Z_57 ;
    wire \generator_inst1.REGSTATZ0Z_58 ;
    wire \generator_inst1.REGSTATZ0Z_59 ;
    wire \generator_inst1.REGSTATZ0Z_53 ;
    wire \generator_inst1.REGSTATZ0Z_54 ;
    wire SELSTAT_c;
    wire \generator_inst1.REGSTATZ0Z_55 ;
    wire \generator_inst1.REGSTATZ0Z_56 ;
    wire _gnd_net_;
    wire CLK_c_g;
    wire SELDYN_c_i_g;
    wire RST_N_c_i_g;

    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__2715),
            .GLOBALBUFFEROUTPUT(CLK_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__2717),
            .DIN(N__2716),
            .DOUT(N__2715),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__2717),
            .PADOUT(N__2716),
            .PADIN(N__2715),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD signal_out_obuf_iopad (
            .OE(N__2706),
            .DIN(N__2705),
            .DOUT(N__2704),
            .PACKAGEPIN(signal_out));
    defparam signal_out_obuf_preio.NEG_TRIGGER=1'b0;
    defparam signal_out_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO signal_out_obuf_preio (
            .PADOEN(N__2706),
            .PADOUT(N__2705),
            .PADIN(N__2704),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1460),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RST_N_ibuf_iopad (
            .OE(N__2697),
            .DIN(N__2696),
            .DOUT(N__2695),
            .PACKAGEPIN(RST_N));
    defparam RST_N_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RST_N_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RST_N_ibuf_preio (
            .PADOEN(N__2697),
            .PADOUT(N__2696),
            .PADIN(N__2695),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RST_N_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SELDYN_ibuf_iopad (
            .OE(N__2688),
            .DIN(N__2687),
            .DOUT(N__2686),
            .PACKAGEPIN(SELDYN));
    defparam SELDYN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SELDYN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SELDYN_ibuf_preio (
            .PADOEN(N__2688),
            .PADOUT(N__2687),
            .PADIN(N__2686),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SELDYN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SELSTAT_ibuf_iopad (
            .OE(N__2679),
            .DIN(N__2678),
            .DOUT(N__2677),
            .PACKAGEPIN(SELSTAT));
    defparam SELSTAT_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SELSTAT_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SELSTAT_ibuf_preio (
            .PADOEN(N__2679),
            .PADOUT(N__2678),
            .PADIN(N__2677),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SELSTAT_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__545 (
            .O(N__2660),
            .I(N__2657));
    LocalMux I__544 (
            .O(N__2657),
            .I(\generator_inst1.REGSTATZ0Z_66 ));
    InMux I__543 (
            .O(N__2654),
            .I(N__2651));
    LocalMux I__542 (
            .O(N__2651),
            .I(\generator_inst1.REGSTATZ0Z_64 ));
    InMux I__541 (
            .O(N__2648),
            .I(N__2645));
    LocalMux I__540 (
            .O(N__2645),
            .I(\generator_inst1.REGSTATZ0Z_65 ));
    InMux I__539 (
            .O(N__2642),
            .I(N__2639));
    LocalMux I__538 (
            .O(N__2639),
            .I(\generator_inst1.REGSTATZ0Z_57 ));
    InMux I__537 (
            .O(N__2636),
            .I(N__2633));
    LocalMux I__536 (
            .O(N__2633),
            .I(\generator_inst1.REGSTATZ0Z_58 ));
    InMux I__535 (
            .O(N__2630),
            .I(N__2627));
    LocalMux I__534 (
            .O(N__2627),
            .I(\generator_inst1.REGSTATZ0Z_59 ));
    InMux I__533 (
            .O(N__2624),
            .I(N__2621));
    LocalMux I__532 (
            .O(N__2621),
            .I(\generator_inst1.REGSTATZ0Z_53 ));
    InMux I__531 (
            .O(N__2618),
            .I(N__2615));
    LocalMux I__530 (
            .O(N__2615),
            .I(\generator_inst1.REGSTATZ0Z_54 ));
    InMux I__529 (
            .O(N__2612),
            .I(N__2560));
    InMux I__528 (
            .O(N__2611),
            .I(N__2560));
    InMux I__527 (
            .O(N__2610),
            .I(N__2549));
    InMux I__526 (
            .O(N__2609),
            .I(N__2549));
    InMux I__525 (
            .O(N__2608),
            .I(N__2549));
    InMux I__524 (
            .O(N__2607),
            .I(N__2549));
    InMux I__523 (
            .O(N__2606),
            .I(N__2549));
    InMux I__522 (
            .O(N__2605),
            .I(N__2540));
    InMux I__521 (
            .O(N__2604),
            .I(N__2540));
    InMux I__520 (
            .O(N__2603),
            .I(N__2540));
    InMux I__519 (
            .O(N__2602),
            .I(N__2540));
    InMux I__518 (
            .O(N__2601),
            .I(N__2515));
    InMux I__517 (
            .O(N__2600),
            .I(N__2515));
    InMux I__516 (
            .O(N__2599),
            .I(N__2515));
    InMux I__515 (
            .O(N__2598),
            .I(N__2515));
    InMux I__514 (
            .O(N__2597),
            .I(N__2515));
    InMux I__513 (
            .O(N__2596),
            .I(N__2500));
    InMux I__512 (
            .O(N__2595),
            .I(N__2500));
    InMux I__511 (
            .O(N__2594),
            .I(N__2500));
    InMux I__510 (
            .O(N__2593),
            .I(N__2500));
    InMux I__509 (
            .O(N__2592),
            .I(N__2500));
    InMux I__508 (
            .O(N__2591),
            .I(N__2500));
    InMux I__507 (
            .O(N__2590),
            .I(N__2500));
    InMux I__506 (
            .O(N__2589),
            .I(N__2491));
    InMux I__505 (
            .O(N__2588),
            .I(N__2491));
    InMux I__504 (
            .O(N__2587),
            .I(N__2491));
    InMux I__503 (
            .O(N__2586),
            .I(N__2491));
    InMux I__502 (
            .O(N__2585),
            .I(N__2476));
    InMux I__501 (
            .O(N__2584),
            .I(N__2476));
    InMux I__500 (
            .O(N__2583),
            .I(N__2476));
    InMux I__499 (
            .O(N__2582),
            .I(N__2476));
    InMux I__498 (
            .O(N__2581),
            .I(N__2476));
    InMux I__497 (
            .O(N__2580),
            .I(N__2476));
    InMux I__496 (
            .O(N__2579),
            .I(N__2476));
    InMux I__495 (
            .O(N__2578),
            .I(N__2459));
    InMux I__494 (
            .O(N__2577),
            .I(N__2459));
    InMux I__493 (
            .O(N__2576),
            .I(N__2459));
    InMux I__492 (
            .O(N__2575),
            .I(N__2459));
    InMux I__491 (
            .O(N__2574),
            .I(N__2459));
    InMux I__490 (
            .O(N__2573),
            .I(N__2459));
    InMux I__489 (
            .O(N__2572),
            .I(N__2459));
    InMux I__488 (
            .O(N__2571),
            .I(N__2459));
    InMux I__487 (
            .O(N__2570),
            .I(N__2446));
    InMux I__486 (
            .O(N__2569),
            .I(N__2446));
    InMux I__485 (
            .O(N__2568),
            .I(N__2446));
    InMux I__484 (
            .O(N__2567),
            .I(N__2446));
    InMux I__483 (
            .O(N__2566),
            .I(N__2446));
    InMux I__482 (
            .O(N__2565),
            .I(N__2446));
    LocalMux I__481 (
            .O(N__2560),
            .I(N__2443));
    LocalMux I__480 (
            .O(N__2549),
            .I(N__2438));
    LocalMux I__479 (
            .O(N__2540),
            .I(N__2438));
    InMux I__478 (
            .O(N__2539),
            .I(N__2425));
    InMux I__477 (
            .O(N__2538),
            .I(N__2425));
    InMux I__476 (
            .O(N__2537),
            .I(N__2425));
    InMux I__475 (
            .O(N__2536),
            .I(N__2425));
    InMux I__474 (
            .O(N__2535),
            .I(N__2425));
    InMux I__473 (
            .O(N__2534),
            .I(N__2425));
    InMux I__472 (
            .O(N__2533),
            .I(N__2408));
    InMux I__471 (
            .O(N__2532),
            .I(N__2408));
    InMux I__470 (
            .O(N__2531),
            .I(N__2408));
    InMux I__469 (
            .O(N__2530),
            .I(N__2408));
    InMux I__468 (
            .O(N__2529),
            .I(N__2408));
    InMux I__467 (
            .O(N__2528),
            .I(N__2408));
    InMux I__466 (
            .O(N__2527),
            .I(N__2408));
    InMux I__465 (
            .O(N__2526),
            .I(N__2408));
    LocalMux I__464 (
            .O(N__2515),
            .I(N__2395));
    LocalMux I__463 (
            .O(N__2500),
            .I(N__2395));
    LocalMux I__462 (
            .O(N__2491),
            .I(N__2395));
    LocalMux I__461 (
            .O(N__2476),
            .I(N__2395));
    LocalMux I__460 (
            .O(N__2459),
            .I(N__2395));
    LocalMux I__459 (
            .O(N__2446),
            .I(N__2395));
    Span4Mux_v I__458 (
            .O(N__2443),
            .I(N__2386));
    Span4Mux_h I__457 (
            .O(N__2438),
            .I(N__2386));
    LocalMux I__456 (
            .O(N__2425),
            .I(N__2386));
    LocalMux I__455 (
            .O(N__2408),
            .I(N__2386));
    Span4Mux_v I__454 (
            .O(N__2395),
            .I(N__2361));
    Span4Mux_v I__453 (
            .O(N__2386),
            .I(N__2358));
    InMux I__452 (
            .O(N__2385),
            .I(N__2345));
    InMux I__451 (
            .O(N__2384),
            .I(N__2345));
    InMux I__450 (
            .O(N__2383),
            .I(N__2345));
    InMux I__449 (
            .O(N__2382),
            .I(N__2345));
    InMux I__448 (
            .O(N__2381),
            .I(N__2345));
    InMux I__447 (
            .O(N__2380),
            .I(N__2345));
    InMux I__446 (
            .O(N__2379),
            .I(N__2328));
    InMux I__445 (
            .O(N__2378),
            .I(N__2328));
    InMux I__444 (
            .O(N__2377),
            .I(N__2328));
    InMux I__443 (
            .O(N__2376),
            .I(N__2328));
    InMux I__442 (
            .O(N__2375),
            .I(N__2328));
    InMux I__441 (
            .O(N__2374),
            .I(N__2328));
    InMux I__440 (
            .O(N__2373),
            .I(N__2328));
    InMux I__439 (
            .O(N__2372),
            .I(N__2328));
    InMux I__438 (
            .O(N__2371),
            .I(N__2305));
    InMux I__437 (
            .O(N__2370),
            .I(N__2305));
    InMux I__436 (
            .O(N__2369),
            .I(N__2305));
    InMux I__435 (
            .O(N__2368),
            .I(N__2305));
    InMux I__434 (
            .O(N__2367),
            .I(N__2305));
    InMux I__433 (
            .O(N__2366),
            .I(N__2305));
    InMux I__432 (
            .O(N__2365),
            .I(N__2305));
    InMux I__431 (
            .O(N__2364),
            .I(N__2305));
    Sp12to4 I__430 (
            .O(N__2361),
            .I(N__2296));
    Sp12to4 I__429 (
            .O(N__2358),
            .I(N__2296));
    LocalMux I__428 (
            .O(N__2345),
            .I(N__2296));
    LocalMux I__427 (
            .O(N__2328),
            .I(N__2296));
    InMux I__426 (
            .O(N__2327),
            .I(N__2283));
    InMux I__425 (
            .O(N__2326),
            .I(N__2283));
    InMux I__424 (
            .O(N__2325),
            .I(N__2283));
    InMux I__423 (
            .O(N__2324),
            .I(N__2283));
    InMux I__422 (
            .O(N__2323),
            .I(N__2283));
    InMux I__421 (
            .O(N__2322),
            .I(N__2283));
    LocalMux I__420 (
            .O(N__2305),
            .I(SELSTAT_c));
    Odrv12 I__419 (
            .O(N__2296),
            .I(SELSTAT_c));
    LocalMux I__418 (
            .O(N__2283),
            .I(SELSTAT_c));
    InMux I__417 (
            .O(N__2276),
            .I(N__2273));
    LocalMux I__416 (
            .O(N__2273),
            .I(\generator_inst1.REGSTATZ0Z_55 ));
    InMux I__415 (
            .O(N__2270),
            .I(N__2267));
    LocalMux I__414 (
            .O(N__2267),
            .I(\generator_inst1.REGSTATZ0Z_56 ));
    ClkMux I__413 (
            .O(N__2264),
            .I(N__2213));
    ClkMux I__412 (
            .O(N__2263),
            .I(N__2213));
    ClkMux I__411 (
            .O(N__2262),
            .I(N__2213));
    ClkMux I__410 (
            .O(N__2261),
            .I(N__2213));
    ClkMux I__409 (
            .O(N__2260),
            .I(N__2213));
    ClkMux I__408 (
            .O(N__2259),
            .I(N__2213));
    ClkMux I__407 (
            .O(N__2258),
            .I(N__2213));
    ClkMux I__406 (
            .O(N__2257),
            .I(N__2213));
    ClkMux I__405 (
            .O(N__2256),
            .I(N__2213));
    ClkMux I__404 (
            .O(N__2255),
            .I(N__2213));
    ClkMux I__403 (
            .O(N__2254),
            .I(N__2213));
    ClkMux I__402 (
            .O(N__2253),
            .I(N__2213));
    ClkMux I__401 (
            .O(N__2252),
            .I(N__2213));
    ClkMux I__400 (
            .O(N__2251),
            .I(N__2213));
    ClkMux I__399 (
            .O(N__2250),
            .I(N__2213));
    ClkMux I__398 (
            .O(N__2249),
            .I(N__2213));
    ClkMux I__397 (
            .O(N__2248),
            .I(N__2213));
    GlobalMux I__396 (
            .O(N__2213),
            .I(N__2210));
    gio2CtrlBuf I__395 (
            .O(N__2210),
            .I(CLK_c_g));
    CEMux I__394 (
            .O(N__2207),
            .I(N__2165));
    CEMux I__393 (
            .O(N__2206),
            .I(N__2165));
    CEMux I__392 (
            .O(N__2205),
            .I(N__2165));
    CEMux I__391 (
            .O(N__2204),
            .I(N__2165));
    CEMux I__390 (
            .O(N__2203),
            .I(N__2165));
    CEMux I__389 (
            .O(N__2202),
            .I(N__2165));
    CEMux I__388 (
            .O(N__2201),
            .I(N__2165));
    CEMux I__387 (
            .O(N__2200),
            .I(N__2165));
    CEMux I__386 (
            .O(N__2199),
            .I(N__2165));
    CEMux I__385 (
            .O(N__2198),
            .I(N__2165));
    CEMux I__384 (
            .O(N__2197),
            .I(N__2165));
    CEMux I__383 (
            .O(N__2196),
            .I(N__2165));
    CEMux I__382 (
            .O(N__2195),
            .I(N__2165));
    CEMux I__381 (
            .O(N__2194),
            .I(N__2165));
    GlobalMux I__380 (
            .O(N__2165),
            .I(N__2162));
    gio2CtrlBuf I__379 (
            .O(N__2162),
            .I(SELDYN_c_i_g));
    SRMux I__378 (
            .O(N__2159),
            .I(N__2108));
    SRMux I__377 (
            .O(N__2158),
            .I(N__2108));
    SRMux I__376 (
            .O(N__2157),
            .I(N__2108));
    SRMux I__375 (
            .O(N__2156),
            .I(N__2108));
    SRMux I__374 (
            .O(N__2155),
            .I(N__2108));
    SRMux I__373 (
            .O(N__2154),
            .I(N__2108));
    SRMux I__372 (
            .O(N__2153),
            .I(N__2108));
    SRMux I__371 (
            .O(N__2152),
            .I(N__2108));
    SRMux I__370 (
            .O(N__2151),
            .I(N__2108));
    SRMux I__369 (
            .O(N__2150),
            .I(N__2108));
    SRMux I__368 (
            .O(N__2149),
            .I(N__2108));
    SRMux I__367 (
            .O(N__2148),
            .I(N__2108));
    SRMux I__366 (
            .O(N__2147),
            .I(N__2108));
    SRMux I__365 (
            .O(N__2146),
            .I(N__2108));
    SRMux I__364 (
            .O(N__2145),
            .I(N__2108));
    SRMux I__363 (
            .O(N__2144),
            .I(N__2108));
    SRMux I__362 (
            .O(N__2143),
            .I(N__2108));
    GlobalMux I__361 (
            .O(N__2108),
            .I(N__2105));
    gio2CtrlBuf I__360 (
            .O(N__2105),
            .I(RST_N_c_i_g));
    InMux I__359 (
            .O(N__2102),
            .I(N__2099));
    LocalMux I__358 (
            .O(N__2099),
            .I(\generator_inst1.REGSTATZ0Z_67 ));
    InMux I__357 (
            .O(N__2096),
            .I(N__2093));
    LocalMux I__356 (
            .O(N__2093),
            .I(\generator_inst1.REGSTATZ0Z_70 ));
    InMux I__355 (
            .O(N__2090),
            .I(N__2087));
    LocalMux I__354 (
            .O(N__2087),
            .I(\generator_inst1.REGSTATZ0Z_68 ));
    InMux I__353 (
            .O(N__2084),
            .I(N__2081));
    LocalMux I__352 (
            .O(N__2081),
            .I(\generator_inst1.REGSTATZ0Z_69 ));
    InMux I__351 (
            .O(N__2078),
            .I(N__2075));
    LocalMux I__350 (
            .O(N__2075),
            .I(\generator_inst1.REGSTATZ0Z_71 ));
    InMux I__349 (
            .O(N__2072),
            .I(N__2069));
    LocalMux I__348 (
            .O(N__2069),
            .I(\generator_inst1.REGSTATZ0Z_72 ));
    InMux I__347 (
            .O(N__2066),
            .I(N__2063));
    LocalMux I__346 (
            .O(N__2063),
            .I(\generator_inst1.REGSTATZ0Z_63 ));
    InMux I__345 (
            .O(N__2060),
            .I(N__2057));
    LocalMux I__344 (
            .O(N__2057),
            .I(\generator_inst1.REGSTATZ0Z_62 ));
    InMux I__343 (
            .O(N__2054),
            .I(N__2051));
    LocalMux I__342 (
            .O(N__2051),
            .I(\generator_inst1.REGSTATZ0Z_60 ));
    InMux I__341 (
            .O(N__2048),
            .I(N__2045));
    LocalMux I__340 (
            .O(N__2045),
            .I(\generator_inst1.REGSTATZ0Z_61 ));
    InMux I__339 (
            .O(N__2042),
            .I(N__2039));
    LocalMux I__338 (
            .O(N__2039),
            .I(\generator_inst1.REGSTATZ0Z_49 ));
    InMux I__337 (
            .O(N__2036),
            .I(N__2033));
    LocalMux I__336 (
            .O(N__2033),
            .I(\generator_inst1.REGSTATZ0Z_50 ));
    InMux I__335 (
            .O(N__2030),
            .I(N__2027));
    LocalMux I__334 (
            .O(N__2027),
            .I(\generator_inst1.REGSTATZ0Z_76 ));
    InMux I__333 (
            .O(N__2024),
            .I(N__2021));
    LocalMux I__332 (
            .O(N__2021),
            .I(\generator_inst1.REGSTATZ0Z_77 ));
    InMux I__331 (
            .O(N__2018),
            .I(N__2015));
    LocalMux I__330 (
            .O(N__2015),
            .I(\generator_inst1.REGSTATZ0Z_78 ));
    InMux I__329 (
            .O(N__2012),
            .I(N__2009));
    LocalMux I__328 (
            .O(N__2009),
            .I(\generator_inst1.REGSTATZ0Z_75 ));
    InMux I__327 (
            .O(N__2006),
            .I(N__2003));
    LocalMux I__326 (
            .O(N__2003),
            .I(\generator_inst1.REGSTATZ0Z_74 ));
    InMux I__325 (
            .O(N__2000),
            .I(N__1997));
    LocalMux I__324 (
            .O(N__1997),
            .I(\generator_inst1.REGSTATZ0Z_73 ));
    InMux I__323 (
            .O(N__1994),
            .I(N__1991));
    LocalMux I__322 (
            .O(N__1991),
            .I(\generator_inst1.REGSTATZ0Z_25 ));
    InMux I__321 (
            .O(N__1988),
            .I(N__1985));
    LocalMux I__320 (
            .O(N__1985),
            .I(\generator_inst1.REGSTATZ0Z_26 ));
    InMux I__319 (
            .O(N__1982),
            .I(N__1979));
    LocalMux I__318 (
            .O(N__1979),
            .I(\generator_inst1.REGSTATZ0Z_30 ));
    InMux I__317 (
            .O(N__1976),
            .I(N__1973));
    LocalMux I__316 (
            .O(N__1973),
            .I(\generator_inst1.REGSTATZ0Z_31 ));
    InMux I__315 (
            .O(N__1970),
            .I(N__1967));
    LocalMux I__314 (
            .O(N__1967),
            .I(\generator_inst1.REGSTATZ0Z_51 ));
    InMux I__313 (
            .O(N__1964),
            .I(N__1961));
    LocalMux I__312 (
            .O(N__1961),
            .I(\generator_inst1.REGSTATZ0Z_52 ));
    InMux I__311 (
            .O(N__1958),
            .I(N__1955));
    LocalMux I__310 (
            .O(N__1955),
            .I(\generator_inst1.REGSTATZ0Z_45 ));
    InMux I__309 (
            .O(N__1952),
            .I(N__1949));
    LocalMux I__308 (
            .O(N__1949),
            .I(\generator_inst1.REGSTATZ0Z_46 ));
    InMux I__307 (
            .O(N__1946),
            .I(N__1943));
    LocalMux I__306 (
            .O(N__1943),
            .I(\generator_inst1.REGSTATZ0Z_47 ));
    InMux I__305 (
            .O(N__1940),
            .I(N__1937));
    LocalMux I__304 (
            .O(N__1937),
            .I(\generator_inst1.REGSTATZ0Z_48 ));
    InMux I__303 (
            .O(N__1934),
            .I(N__1931));
    LocalMux I__302 (
            .O(N__1931),
            .I(\generator_inst1.REGSTATZ0Z_19 ));
    InMux I__301 (
            .O(N__1928),
            .I(N__1925));
    LocalMux I__300 (
            .O(N__1925),
            .I(\generator_inst1.REGSTATZ0Z_22 ));
    InMux I__299 (
            .O(N__1922),
            .I(N__1919));
    LocalMux I__298 (
            .O(N__1919),
            .I(\generator_inst1.REGSTATZ0Z_20 ));
    InMux I__297 (
            .O(N__1916),
            .I(N__1913));
    LocalMux I__296 (
            .O(N__1913),
            .I(\generator_inst1.REGSTATZ0Z_21 ));
    InMux I__295 (
            .O(N__1910),
            .I(N__1907));
    LocalMux I__294 (
            .O(N__1907),
            .I(\generator_inst1.REGSTATZ0Z_0 ));
    InMux I__293 (
            .O(N__1904),
            .I(N__1901));
    LocalMux I__292 (
            .O(N__1901),
            .I(\generator_inst1.REGSTATZ0Z_1 ));
    InMux I__291 (
            .O(N__1898),
            .I(N__1895));
    LocalMux I__290 (
            .O(N__1895),
            .I(\generator_inst1.REGSTATZ0Z_27 ));
    InMux I__289 (
            .O(N__1892),
            .I(N__1889));
    LocalMux I__288 (
            .O(N__1889),
            .I(\generator_inst1.REGSTATZ0Z_28 ));
    InMux I__287 (
            .O(N__1886),
            .I(N__1883));
    LocalMux I__286 (
            .O(N__1883),
            .I(\generator_inst1.REGSTATZ0Z_29 ));
    InMux I__285 (
            .O(N__1880),
            .I(N__1877));
    LocalMux I__284 (
            .O(N__1877),
            .I(\generator_inst1.REGSTATZ0Z_79 ));
    InMux I__283 (
            .O(N__1874),
            .I(N__1871));
    LocalMux I__282 (
            .O(N__1871),
            .I(\generator_inst1.REGSTATZ0Z_82 ));
    InMux I__281 (
            .O(N__1868),
            .I(N__1865));
    LocalMux I__280 (
            .O(N__1865),
            .I(\generator_inst1.REGSTATZ0Z_83 ));
    InMux I__279 (
            .O(N__1862),
            .I(N__1859));
    LocalMux I__278 (
            .O(N__1859),
            .I(\generator_inst1.REGSTATZ0Z_5 ));
    InMux I__277 (
            .O(N__1856),
            .I(N__1853));
    LocalMux I__276 (
            .O(N__1853),
            .I(\generator_inst1.REGSTATZ0Z_2 ));
    InMux I__275 (
            .O(N__1850),
            .I(N__1847));
    LocalMux I__274 (
            .O(N__1847),
            .I(\generator_inst1.REGSTATZ0Z_3 ));
    InMux I__273 (
            .O(N__1844),
            .I(N__1841));
    LocalMux I__272 (
            .O(N__1841),
            .I(\generator_inst1.REGSTATZ0Z_4 ));
    InMux I__271 (
            .O(N__1838),
            .I(N__1835));
    LocalMux I__270 (
            .O(N__1835),
            .I(\generator_inst1.REGSTATZ0Z_24 ));
    InMux I__269 (
            .O(N__1832),
            .I(N__1829));
    LocalMux I__268 (
            .O(N__1829),
            .I(\generator_inst1.REGSTATZ0Z_23 ));
    InMux I__267 (
            .O(N__1826),
            .I(N__1823));
    LocalMux I__266 (
            .O(N__1823),
            .I(\generator_inst1.REGSTATZ0Z_40 ));
    InMux I__265 (
            .O(N__1820),
            .I(N__1817));
    LocalMux I__264 (
            .O(N__1817),
            .I(\generator_inst1.REGSTATZ0Z_41 ));
    InMux I__263 (
            .O(N__1814),
            .I(N__1811));
    LocalMux I__262 (
            .O(N__1811),
            .I(\generator_inst1.REGSTATZ0Z_42 ));
    InMux I__261 (
            .O(N__1808),
            .I(N__1805));
    LocalMux I__260 (
            .O(N__1805),
            .I(\generator_inst1.REGSTATZ0Z_43 ));
    InMux I__259 (
            .O(N__1802),
            .I(N__1799));
    LocalMux I__258 (
            .O(N__1799),
            .I(\generator_inst1.REGSTATZ0Z_44 ));
    InMux I__257 (
            .O(N__1796),
            .I(N__1793));
    LocalMux I__256 (
            .O(N__1793),
            .I(N__1790));
    Span4Mux_v I__255 (
            .O(N__1790),
            .I(N__1769));
    InMux I__254 (
            .O(N__1789),
            .I(N__1764));
    InMux I__253 (
            .O(N__1788),
            .I(N__1764));
    InMux I__252 (
            .O(N__1787),
            .I(N__1747));
    InMux I__251 (
            .O(N__1786),
            .I(N__1747));
    InMux I__250 (
            .O(N__1785),
            .I(N__1747));
    InMux I__249 (
            .O(N__1784),
            .I(N__1747));
    InMux I__248 (
            .O(N__1783),
            .I(N__1747));
    InMux I__247 (
            .O(N__1782),
            .I(N__1747));
    InMux I__246 (
            .O(N__1781),
            .I(N__1747));
    InMux I__245 (
            .O(N__1780),
            .I(N__1747));
    InMux I__244 (
            .O(N__1779),
            .I(N__1730));
    InMux I__243 (
            .O(N__1778),
            .I(N__1730));
    InMux I__242 (
            .O(N__1777),
            .I(N__1730));
    InMux I__241 (
            .O(N__1776),
            .I(N__1730));
    InMux I__240 (
            .O(N__1775),
            .I(N__1730));
    InMux I__239 (
            .O(N__1774),
            .I(N__1730));
    InMux I__238 (
            .O(N__1773),
            .I(N__1730));
    InMux I__237 (
            .O(N__1772),
            .I(N__1730));
    Span4Mux_v I__236 (
            .O(N__1769),
            .I(N__1721));
    LocalMux I__235 (
            .O(N__1764),
            .I(N__1721));
    LocalMux I__234 (
            .O(N__1747),
            .I(N__1721));
    LocalMux I__233 (
            .O(N__1730),
            .I(N__1721));
    Span4Mux_v I__232 (
            .O(N__1721),
            .I(N__1718));
    Span4Mux_v I__231 (
            .O(N__1718),
            .I(N__1715));
    Odrv4 I__230 (
            .O(N__1715),
            .I(SELDYN_c));
    IoInMux I__229 (
            .O(N__1712),
            .I(N__1709));
    LocalMux I__228 (
            .O(N__1709),
            .I(SELDYN_c_i));
    InMux I__227 (
            .O(N__1706),
            .I(N__1703));
    LocalMux I__226 (
            .O(N__1703),
            .I(N__1700));
    Span4Mux_v I__225 (
            .O(N__1700),
            .I(N__1697));
    Span4Mux_v I__224 (
            .O(N__1697),
            .I(N__1694));
    Odrv4 I__223 (
            .O(N__1694),
            .I(RST_N_c));
    IoInMux I__222 (
            .O(N__1691),
            .I(N__1688));
    LocalMux I__221 (
            .O(N__1688),
            .I(N__1685));
    IoSpan4Mux I__220 (
            .O(N__1685),
            .I(N__1682));
    Odrv4 I__219 (
            .O(N__1682),
            .I(RST_N_c_i));
    InMux I__218 (
            .O(N__1679),
            .I(N__1676));
    LocalMux I__217 (
            .O(N__1676),
            .I(\generator_inst1.REGSTATZ0Z_80 ));
    InMux I__216 (
            .O(N__1673),
            .I(N__1670));
    LocalMux I__215 (
            .O(N__1670),
            .I(\generator_inst1.REGSTATZ0Z_81 ));
    InMux I__214 (
            .O(N__1667),
            .I(N__1664));
    LocalMux I__213 (
            .O(N__1664),
            .I(\generator_inst1.REGSTATZ0Z_34 ));
    InMux I__212 (
            .O(N__1661),
            .I(N__1658));
    LocalMux I__211 (
            .O(N__1658),
            .I(\generator_inst1.REGSTATZ0Z_35 ));
    InMux I__210 (
            .O(N__1655),
            .I(N__1652));
    LocalMux I__209 (
            .O(N__1652),
            .I(\generator_inst1.REGSTATZ0Z_36 ));
    InMux I__208 (
            .O(N__1649),
            .I(N__1646));
    LocalMux I__207 (
            .O(N__1646),
            .I(\generator_inst1.REGSTATZ0Z_32 ));
    InMux I__206 (
            .O(N__1643),
            .I(N__1640));
    LocalMux I__205 (
            .O(N__1640),
            .I(\generator_inst1.REGSTATZ0Z_33 ));
    InMux I__204 (
            .O(N__1637),
            .I(N__1634));
    LocalMux I__203 (
            .O(N__1634),
            .I(\generator_inst1.REGSTATZ0Z_37 ));
    InMux I__202 (
            .O(N__1631),
            .I(N__1628));
    LocalMux I__201 (
            .O(N__1628),
            .I(\generator_inst1.REGSTATZ0Z_38 ));
    InMux I__200 (
            .O(N__1625),
            .I(N__1622));
    LocalMux I__199 (
            .O(N__1622),
            .I(\generator_inst1.REGSTATZ0Z_39 ));
    InMux I__198 (
            .O(N__1619),
            .I(N__1616));
    LocalMux I__197 (
            .O(N__1616),
            .I(\generator_inst1.REGSTATZ0Z_10 ));
    InMux I__196 (
            .O(N__1613),
            .I(N__1610));
    LocalMux I__195 (
            .O(N__1610),
            .I(\generator_inst1.REGSTATZ0Z_11 ));
    InMux I__194 (
            .O(N__1607),
            .I(N__1604));
    LocalMux I__193 (
            .O(N__1604),
            .I(\generator_inst1.REGSTATZ0Z_12 ));
    InMux I__192 (
            .O(N__1601),
            .I(N__1598));
    LocalMux I__191 (
            .O(N__1598),
            .I(\generator_inst1.REGSTATZ0Z_13 ));
    InMux I__190 (
            .O(N__1595),
            .I(N__1592));
    LocalMux I__189 (
            .O(N__1592),
            .I(\generator_inst1.REGSTATZ0Z_18 ));
    InMux I__188 (
            .O(N__1589),
            .I(N__1586));
    LocalMux I__187 (
            .O(N__1586),
            .I(\generator_inst1.REGSTATZ0Z_14 ));
    InMux I__186 (
            .O(N__1583),
            .I(N__1580));
    LocalMux I__185 (
            .O(N__1580),
            .I(\generator_inst1.REGSTATZ0Z_15 ));
    InMux I__184 (
            .O(N__1577),
            .I(N__1574));
    LocalMux I__183 (
            .O(N__1574),
            .I(\generator_inst1.REGSTATZ0Z_16 ));
    InMux I__182 (
            .O(N__1571),
            .I(N__1568));
    LocalMux I__181 (
            .O(N__1568),
            .I(\generator_inst1.REGSTATZ0Z_17 ));
    InMux I__180 (
            .O(N__1565),
            .I(N__1562));
    LocalMux I__179 (
            .O(N__1562),
            .I(\generator_inst1.REGSTATZ0Z_86 ));
    CascadeMux I__178 (
            .O(N__1559),
            .I(N__1556));
    InMux I__177 (
            .O(N__1556),
            .I(N__1553));
    LocalMux I__176 (
            .O(N__1553),
            .I(\generator_inst1.REGSTATZ0Z_87 ));
    InMux I__175 (
            .O(N__1550),
            .I(N__1547));
    LocalMux I__174 (
            .O(N__1547),
            .I(\generator_inst1.REGSTATZ0Z_84 ));
    InMux I__173 (
            .O(N__1544),
            .I(N__1541));
    LocalMux I__172 (
            .O(N__1541),
            .I(\generator_inst1.REGSTATZ0Z_85 ));
    InMux I__171 (
            .O(N__1538),
            .I(N__1535));
    LocalMux I__170 (
            .O(N__1535),
            .I(\generator_inst1.REGSTATZ0Z_9 ));
    InMux I__169 (
            .O(N__1532),
            .I(N__1529));
    LocalMux I__168 (
            .O(N__1529),
            .I(\generator_inst1.REGSTATZ0Z_6 ));
    InMux I__167 (
            .O(N__1526),
            .I(N__1523));
    LocalMux I__166 (
            .O(N__1523),
            .I(\generator_inst1.REGSTATZ0Z_7 ));
    InMux I__165 (
            .O(N__1520),
            .I(N__1517));
    LocalMux I__164 (
            .O(N__1517),
            .I(\generator_inst1.REGSTATZ0Z_8 ));
    InMux I__163 (
            .O(N__1514),
            .I(N__1511));
    LocalMux I__162 (
            .O(N__1511),
            .I(\generator_inst1.REGDYNZ0Z_11 ));
    InMux I__161 (
            .O(N__1508),
            .I(N__1505));
    LocalMux I__160 (
            .O(N__1505),
            .I(\generator_inst1.REGDYNZ0Z_12 ));
    InMux I__159 (
            .O(N__1502),
            .I(N__1499));
    LocalMux I__158 (
            .O(N__1499),
            .I(\generator_inst1.REGDYNZ0Z_13 ));
    InMux I__157 (
            .O(N__1496),
            .I(N__1493));
    LocalMux I__156 (
            .O(N__1493),
            .I(\generator_inst1.REGDYNZ0Z_14 ));
    InMux I__155 (
            .O(N__1490),
            .I(N__1487));
    LocalMux I__154 (
            .O(N__1487),
            .I(\generator_inst1.REGDYNZ0Z_9 ));
    InMux I__153 (
            .O(N__1484),
            .I(N__1481));
    LocalMux I__152 (
            .O(N__1481),
            .I(\generator_inst1.REGDYNZ0Z_7 ));
    InMux I__151 (
            .O(N__1478),
            .I(N__1475));
    LocalMux I__150 (
            .O(N__1475),
            .I(\generator_inst1.REGDYNZ0Z_8 ));
    InMux I__149 (
            .O(N__1472),
            .I(N__1469));
    LocalMux I__148 (
            .O(N__1469),
            .I(\generator_inst1.REGDYNZ0Z_15 ));
    InMux I__147 (
            .O(N__1466),
            .I(N__1463));
    LocalMux I__146 (
            .O(N__1463),
            .I(generated_signal));
    IoInMux I__145 (
            .O(N__1460),
            .I(N__1457));
    LocalMux I__144 (
            .O(N__1457),
            .I(N__1454));
    Span4Mux_s1_h I__143 (
            .O(N__1454),
            .I(N__1451));
    Span4Mux_v I__142 (
            .O(N__1451),
            .I(N__1448));
    Odrv4 I__141 (
            .O(N__1448),
            .I(signal_out_c));
    CEMux I__140 (
            .O(N__1445),
            .I(N__1442));
    LocalMux I__139 (
            .O(N__1442),
            .I(N__1439));
    Sp12to4 I__138 (
            .O(N__1439),
            .I(N__1435));
    CEMux I__137 (
            .O(N__1438),
            .I(N__1432));
    Odrv12 I__136 (
            .O(N__1435),
            .I(\generator_inst1.REGDYN8_iZ0 ));
    LocalMux I__135 (
            .O(N__1432),
            .I(\generator_inst1.REGDYN8_iZ0 ));
    InMux I__134 (
            .O(N__1427),
            .I(N__1424));
    LocalMux I__133 (
            .O(N__1424),
            .I(\generator_inst1.REGDYNZ0Z_1 ));
    InMux I__132 (
            .O(N__1421),
            .I(N__1418));
    LocalMux I__131 (
            .O(N__1418),
            .I(\generator_inst1.REGDYNZ0Z_2 ));
    InMux I__130 (
            .O(N__1415),
            .I(N__1412));
    LocalMux I__129 (
            .O(N__1412),
            .I(\generator_inst1.REGDYNZ0Z_5 ));
    InMux I__128 (
            .O(N__1409),
            .I(N__1406));
    LocalMux I__127 (
            .O(N__1406),
            .I(\generator_inst1.REGDYNZ0Z_6 ));
    InMux I__126 (
            .O(N__1403),
            .I(N__1400));
    LocalMux I__125 (
            .O(N__1400),
            .I(\generator_inst1.REGDYNZ0Z_3 ));
    InMux I__124 (
            .O(N__1397),
            .I(N__1394));
    LocalMux I__123 (
            .O(N__1394),
            .I(\generator_inst1.REGDYNZ0Z_4 ));
    InMux I__122 (
            .O(N__1391),
            .I(N__1388));
    LocalMux I__121 (
            .O(N__1388),
            .I(\generator_inst1.REGDYNZ0Z_0 ));
    InMux I__120 (
            .O(N__1385),
            .I(N__1382));
    LocalMux I__119 (
            .O(N__1382),
            .I(\generator_inst1.REGDYNZ0Z_10 ));
    ICE_GB RST_N_ibuf_RNIBJGC_0 (
            .USERSIGNALTOGLOBALBUFFER(N__1691),
            .GLOBALBUFFEROUTPUT(RST_N_c_i_g));
    GND GND (
            .Y(GNDG0));
    ICE_GB SELDYN_ibuf_RNIKHL3_0 (
            .USERSIGNALTOGLOBALBUFFER(N__1712),
            .GLOBALBUFFEROUTPUT(SELDYN_c_i_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \generator_inst1.REGDYN_2_LC_1_9_0 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_2_LC_1_9_0 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_2_LC_1_9_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGDYN_2_LC_1_9_0  (
            .in0(N__1774),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1427),
            .lcout(\generator_inst1.REGDYNZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2264),
            .ce(N__1445),
            .sr(N__2159));
    defparam \generator_inst1.REGDYN_1_LC_1_9_1 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_1_LC_1_9_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGDYN_1_LC_1_9_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGDYN_1_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(N__1773),
            .in2(_gnd_net_),
            .in3(N__1391),
            .lcout(\generator_inst1.REGDYNZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2264),
            .ce(N__1445),
            .sr(N__2159));
    defparam \generator_inst1.REGDYN_3_LC_1_9_2 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_3_LC_1_9_2 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_3_LC_1_9_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGDYN_3_LC_1_9_2  (
            .in0(N__1775),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1421),
            .lcout(\generator_inst1.REGDYNZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2264),
            .ce(N__1445),
            .sr(N__2159));
    defparam \generator_inst1.REGDYN_7_LC_1_9_3 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_7_LC_1_9_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_7_LC_1_9_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGDYN_7_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(N__1779),
            .in2(_gnd_net_),
            .in3(N__1409),
            .lcout(\generator_inst1.REGDYNZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2264),
            .ce(N__1445),
            .sr(N__2159));
    defparam \generator_inst1.REGDYN_5_LC_1_9_4 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_5_LC_1_9_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGDYN_5_LC_1_9_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGDYN_5_LC_1_9_4  (
            .in0(N__1777),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1397),
            .lcout(\generator_inst1.REGDYNZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2264),
            .ce(N__1445),
            .sr(N__2159));
    defparam \generator_inst1.REGDYN_6_LC_1_9_5 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_6_LC_1_9_5 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_6_LC_1_9_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGDYN_6_LC_1_9_5  (
            .in0(_gnd_net_),
            .in1(N__1778),
            .in2(_gnd_net_),
            .in3(N__1415),
            .lcout(\generator_inst1.REGDYNZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2264),
            .ce(N__1445),
            .sr(N__2159));
    defparam \generator_inst1.REGDYN_4_LC_1_9_6 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_4_LC_1_9_6 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGDYN_4_LC_1_9_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGDYN_4_LC_1_9_6  (
            .in0(N__1776),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1403),
            .lcout(\generator_inst1.REGDYNZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2264),
            .ce(N__1445),
            .sr(N__2159));
    defparam \generator_inst1.REGDYN_0_LC_1_9_7 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_0_LC_1_9_7 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_0_LC_1_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \generator_inst1.REGDYN_0_LC_1_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1772),
            .lcout(\generator_inst1.REGDYNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2264),
            .ce(N__1445),
            .sr(N__2159));
    defparam \generator_inst1.REGDYN_11_LC_1_10_0 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_11_LC_1_10_0 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_11_LC_1_10_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGDYN_11_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__1781),
            .in2(_gnd_net_),
            .in3(N__1385),
            .lcout(\generator_inst1.REGDYNZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2263),
            .ce(N__1438),
            .sr(N__2158));
    defparam \generator_inst1.REGDYN_10_LC_1_10_1 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_10_LC_1_10_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGDYN_10_LC_1_10_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGDYN_10_LC_1_10_1  (
            .in0(N__1780),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1490),
            .lcout(\generator_inst1.REGDYNZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2263),
            .ce(N__1438),
            .sr(N__2158));
    defparam \generator_inst1.REGDYN_12_LC_1_10_2 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_12_LC_1_10_2 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGDYN_12_LC_1_10_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGDYN_12_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__1782),
            .in2(_gnd_net_),
            .in3(N__1514),
            .lcout(\generator_inst1.REGDYNZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2263),
            .ce(N__1438),
            .sr(N__2158));
    defparam \generator_inst1.REGDYN_13_LC_1_10_3 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_13_LC_1_10_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_13_LC_1_10_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGDYN_13_LC_1_10_3  (
            .in0(N__1783),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1508),
            .lcout(\generator_inst1.REGDYNZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2263),
            .ce(N__1438),
            .sr(N__2158));
    defparam \generator_inst1.REGDYN_14_LC_1_10_4 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_14_LC_1_10_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGDYN_14_LC_1_10_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGDYN_14_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(N__1784),
            .in2(_gnd_net_),
            .in3(N__1502),
            .lcout(\generator_inst1.REGDYNZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2263),
            .ce(N__1438),
            .sr(N__2158));
    defparam \generator_inst1.REGDYN_15_LC_1_10_5 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_15_LC_1_10_5 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_15_LC_1_10_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGDYN_15_LC_1_10_5  (
            .in0(N__1785),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1496),
            .lcout(\generator_inst1.REGDYNZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2263),
            .ce(N__1438),
            .sr(N__2158));
    defparam \generator_inst1.REGDYN_9_LC_1_10_6 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_9_LC_1_10_6 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_9_LC_1_10_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGDYN_9_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(N__1787),
            .in2(_gnd_net_),
            .in3(N__1478),
            .lcout(\generator_inst1.REGDYNZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2263),
            .ce(N__1438),
            .sr(N__2158));
    defparam \generator_inst1.REGDYN_8_LC_1_10_7 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_8_LC_1_10_7 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_8_LC_1_10_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGDYN_8_LC_1_10_7  (
            .in0(N__1786),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1484),
            .lcout(\generator_inst1.REGDYNZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2263),
            .ce(N__1438),
            .sr(N__2158));
    defparam \generator_inst1.signal_out_LC_1_11_0 .C_ON=1'b0;
    defparam \generator_inst1.signal_out_LC_1_11_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.signal_out_LC_1_11_0 .LUT_INIT=16'b0110001001000000;
    LogicCell40 \generator_inst1.signal_out_LC_1_11_0  (
            .in0(N__2612),
            .in1(N__1789),
            .in2(N__1559),
            .in3(N__1472),
            .lcout(generated_signal),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2260),
            .ce(),
            .sr(N__2155));
    defparam \receptor_inst1.signal_out_LC_1_11_1 .C_ON=1'b0;
    defparam \receptor_inst1.signal_out_LC_1_11_1 .SEQ_MODE=4'b1010;
    defparam \receptor_inst1.signal_out_LC_1_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \receptor_inst1.signal_out_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1466),
            .lcout(signal_out_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2260),
            .ce(),
            .sr(N__2155));
    defparam \generator_inst1.REGDYN8_i_LC_1_11_2 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN8_i_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.REGDYN8_i_LC_1_11_2 .LUT_INIT=16'b1101110111011101;
    LogicCell40 \generator_inst1.REGDYN8_i_LC_1_11_2  (
            .in0(N__2611),
            .in1(N__1788),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\generator_inst1.REGDYN8_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.REGSTAT_86_LC_1_12_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_86_LC_1_12_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_86_LC_1_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_86_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__2604),
            .in2(_gnd_net_),
            .in3(N__1544),
            .lcout(\generator_inst1.REGSTATZ0Z_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2257),
            .ce(N__2203),
            .sr(N__2152));
    defparam \generator_inst1.REGSTAT_87_LC_1_12_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_87_LC_1_12_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_87_LC_1_12_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_87_LC_1_12_1  (
            .in0(N__2605),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1565),
            .lcout(\generator_inst1.REGSTATZ0Z_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2257),
            .ce(N__2203),
            .sr(N__2152));
    defparam \generator_inst1.REGSTAT_84_LC_1_12_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_84_LC_1_12_5 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_84_LC_1_12_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_84_LC_1_12_5  (
            .in0(N__2602),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1868),
            .lcout(\generator_inst1.REGSTATZ0Z_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2257),
            .ce(N__2203),
            .sr(N__2152));
    defparam \generator_inst1.REGSTAT_85_LC_1_12_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_85_LC_1_12_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_85_LC_1_12_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_85_LC_1_12_7  (
            .in0(N__2603),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1550),
            .lcout(\generator_inst1.REGSTATZ0Z_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2257),
            .ce(N__2203),
            .sr(N__2152));
    defparam \generator_inst1.REGSTAT_10_LC_1_13_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_10_LC_1_13_0 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_10_LC_1_13_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_10_LC_1_13_0  (
            .in0(N__2534),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1538),
            .lcout(\generator_inst1.REGSTATZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2254),
            .ce(N__2200),
            .sr(N__2149));
    defparam \generator_inst1.REGSTAT_7_LC_1_13_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_7_LC_1_13_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_7_LC_1_13_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_7_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__2537),
            .in2(_gnd_net_),
            .in3(N__1532),
            .lcout(\generator_inst1.REGSTATZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2254),
            .ce(N__2200),
            .sr(N__2149));
    defparam \generator_inst1.REGSTAT_9_LC_1_13_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_9_LC_1_13_2 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_9_LC_1_13_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_9_LC_1_13_2  (
            .in0(N__2539),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1520),
            .lcout(\generator_inst1.REGSTATZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2254),
            .ce(N__2200),
            .sr(N__2149));
    defparam \generator_inst1.REGSTAT_6_LC_1_13_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_6_LC_1_13_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_6_LC_1_13_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_6_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__2536),
            .in2(_gnd_net_),
            .in3(N__1862),
            .lcout(\generator_inst1.REGSTATZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2254),
            .ce(N__2200),
            .sr(N__2149));
    defparam \generator_inst1.REGSTAT_8_LC_1_13_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_8_LC_1_13_5 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_8_LC_1_13_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_8_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__2538),
            .in2(_gnd_net_),
            .in3(N__1526),
            .lcout(\generator_inst1.REGSTATZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2254),
            .ce(N__2200),
            .sr(N__2149));
    defparam \generator_inst1.REGSTAT_11_LC_1_13_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_11_LC_1_13_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_11_LC_1_13_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_11_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__2535),
            .in2(_gnd_net_),
            .in3(N__1619),
            .lcout(\generator_inst1.REGSTATZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2254),
            .ce(N__2200),
            .sr(N__2149));
    defparam \generator_inst1.REGSTAT_19_LC_1_14_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_19_LC_1_14_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_19_LC_1_14_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_19_LC_1_14_0  (
            .in0(N__2533),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1595),
            .lcout(\generator_inst1.REGSTATZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2251),
            .ce(N__2197),
            .sr(N__2147));
    defparam \generator_inst1.REGSTAT_12_LC_1_14_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_12_LC_1_14_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_12_LC_1_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_12_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__2526),
            .in2(_gnd_net_),
            .in3(N__1613),
            .lcout(\generator_inst1.REGSTATZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2251),
            .ce(N__2197),
            .sr(N__2147));
    defparam \generator_inst1.REGSTAT_14_LC_1_14_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_14_LC_1_14_2 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_14_LC_1_14_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_14_LC_1_14_2  (
            .in0(N__2528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1601),
            .lcout(\generator_inst1.REGSTATZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2251),
            .ce(N__2197),
            .sr(N__2147));
    defparam \generator_inst1.REGSTAT_13_LC_1_14_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_13_LC_1_14_3 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_13_LC_1_14_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_13_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__2527),
            .in2(_gnd_net_),
            .in3(N__1607),
            .lcout(\generator_inst1.REGSTATZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2251),
            .ce(N__2197),
            .sr(N__2147));
    defparam \generator_inst1.REGSTAT_18_LC_1_14_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_18_LC_1_14_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_18_LC_1_14_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_18_LC_1_14_4  (
            .in0(N__2532),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1571),
            .lcout(\generator_inst1.REGSTATZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2251),
            .ce(N__2197),
            .sr(N__2147));
    defparam \generator_inst1.REGSTAT_15_LC_1_14_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_15_LC_1_14_5 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_15_LC_1_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_15_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__2529),
            .in2(_gnd_net_),
            .in3(N__1589),
            .lcout(\generator_inst1.REGSTATZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2251),
            .ce(N__2197),
            .sr(N__2147));
    defparam \generator_inst1.REGSTAT_16_LC_1_14_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_16_LC_1_14_6 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_16_LC_1_14_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_16_LC_1_14_6  (
            .in0(N__2530),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1583),
            .lcout(\generator_inst1.REGSTATZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2251),
            .ce(N__2197),
            .sr(N__2147));
    defparam \generator_inst1.REGSTAT_17_LC_1_14_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_17_LC_1_14_7 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_17_LC_1_14_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_17_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(N__2531),
            .in2(_gnd_net_),
            .in3(N__1577),
            .lcout(\generator_inst1.REGSTATZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2251),
            .ce(N__2197),
            .sr(N__2147));
    defparam \generator_inst1.REGSTAT_32_LC_1_15_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_32_LC_1_15_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_32_LC_1_15_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_32_LC_1_15_0  (
            .in0(N__2364),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1976),
            .lcout(\generator_inst1.REGSTATZ0Z_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2249),
            .ce(N__2195),
            .sr(N__2145));
    defparam \generator_inst1.REGSTAT_34_LC_1_15_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_34_LC_1_15_1 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_34_LC_1_15_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_34_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__2366),
            .in2(_gnd_net_),
            .in3(N__1643),
            .lcout(\generator_inst1.REGSTATZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2249),
            .ce(N__2195),
            .sr(N__2145));
    defparam \generator_inst1.REGSTAT_37_LC_1_15_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_37_LC_1_15_2 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_37_LC_1_15_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_37_LC_1_15_2  (
            .in0(N__2369),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1655),
            .lcout(\generator_inst1.REGSTATZ0Z_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2249),
            .ce(N__2195),
            .sr(N__2145));
    defparam \generator_inst1.REGSTAT_35_LC_1_15_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_35_LC_1_15_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_35_LC_1_15_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_35_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__2367),
            .in2(_gnd_net_),
            .in3(N__1667),
            .lcout(\generator_inst1.REGSTATZ0Z_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2249),
            .ce(N__2195),
            .sr(N__2145));
    defparam \generator_inst1.REGSTAT_36_LC_1_15_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_36_LC_1_15_4 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_36_LC_1_15_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_36_LC_1_15_4  (
            .in0(N__2368),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1661),
            .lcout(\generator_inst1.REGSTATZ0Z_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2249),
            .ce(N__2195),
            .sr(N__2145));
    defparam \generator_inst1.REGSTAT_39_LC_1_15_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_39_LC_1_15_5 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_39_LC_1_15_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_39_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__2371),
            .in2(_gnd_net_),
            .in3(N__1631),
            .lcout(\generator_inst1.REGSTATZ0Z_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2249),
            .ce(N__2195),
            .sr(N__2145));
    defparam \generator_inst1.REGSTAT_33_LC_1_15_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_33_LC_1_15_6 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_33_LC_1_15_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_33_LC_1_15_6  (
            .in0(N__2365),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1649),
            .lcout(\generator_inst1.REGSTATZ0Z_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2249),
            .ce(N__2195),
            .sr(N__2145));
    defparam \generator_inst1.REGSTAT_38_LC_1_15_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_38_LC_1_15_7 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_38_LC_1_15_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_38_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(N__2370),
            .in2(_gnd_net_),
            .in3(N__1637),
            .lcout(\generator_inst1.REGSTATZ0Z_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2249),
            .ce(N__2195),
            .sr(N__2145));
    defparam \generator_inst1.REGSTAT_41_LC_1_16_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_41_LC_1_16_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_41_LC_1_16_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_41_LC_1_16_0  (
            .in0(N__2323),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1826),
            .lcout(\generator_inst1.REGSTATZ0Z_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2248),
            .ce(N__2194),
            .sr(N__2143));
    defparam \generator_inst1.REGSTAT_40_LC_1_16_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_40_LC_1_16_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_40_LC_1_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_40_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(N__2322),
            .in2(_gnd_net_),
            .in3(N__1625),
            .lcout(\generator_inst1.REGSTATZ0Z_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2248),
            .ce(N__2194),
            .sr(N__2143));
    defparam \generator_inst1.REGSTAT_44_LC_1_16_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_44_LC_1_16_2 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_44_LC_1_16_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_44_LC_1_16_2  (
            .in0(N__2326),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1808),
            .lcout(\generator_inst1.REGSTATZ0Z_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2248),
            .ce(N__2194),
            .sr(N__2143));
    defparam \generator_inst1.REGSTAT_42_LC_1_16_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_42_LC_1_16_4 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_42_LC_1_16_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_42_LC_1_16_4  (
            .in0(N__2324),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1820),
            .lcout(\generator_inst1.REGSTATZ0Z_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2248),
            .ce(N__2194),
            .sr(N__2143));
    defparam \generator_inst1.REGSTAT_43_LC_1_16_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_43_LC_1_16_5 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_43_LC_1_16_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_43_LC_1_16_5  (
            .in0(_gnd_net_),
            .in1(N__2325),
            .in2(_gnd_net_),
            .in3(N__1814),
            .lcout(\generator_inst1.REGSTATZ0Z_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2248),
            .ce(N__2194),
            .sr(N__2143));
    defparam \generator_inst1.REGSTAT_45_LC_1_16_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_45_LC_1_16_6 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_45_LC_1_16_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_45_LC_1_16_6  (
            .in0(N__2327),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1802),
            .lcout(\generator_inst1.REGSTATZ0Z_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2248),
            .ce(N__2194),
            .sr(N__2143));
    defparam SELDYN_ibuf_RNIKHL3_LC_1_17_3.C_ON=1'b0;
    defparam SELDYN_ibuf_RNIKHL3_LC_1_17_3.SEQ_MODE=4'b0000;
    defparam SELDYN_ibuf_RNIKHL3_LC_1_17_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 SELDYN_ibuf_RNIKHL3_LC_1_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1796),
            .lcout(SELDYN_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RST_N_ibuf_RNIBJGC_LC_1_18_5.C_ON=1'b0;
    defparam RST_N_ibuf_RNIBJGC_LC_1_18_5.SEQ_MODE=4'b0000;
    defparam RST_N_ibuf_RNIBJGC_LC_1_18_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 RST_N_ibuf_RNIBJGC_LC_1_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1706),
            .lcout(RST_N_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.REGSTAT_80_LC_2_12_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_80_LC_2_12_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_80_LC_2_12_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_80_LC_2_12_0  (
            .in0(N__2607),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1880),
            .lcout(\generator_inst1.REGSTATZ0Z_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2261),
            .ce(N__2206),
            .sr(N__2156));
    defparam \generator_inst1.REGSTAT_82_LC_2_12_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_82_LC_2_12_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_82_LC_2_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_82_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__2609),
            .in2(_gnd_net_),
            .in3(N__1673),
            .lcout(\generator_inst1.REGSTATZ0Z_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2261),
            .ce(N__2206),
            .sr(N__2156));
    defparam \generator_inst1.REGSTAT_81_LC_2_12_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_81_LC_2_12_2 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_81_LC_2_12_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_81_LC_2_12_2  (
            .in0(N__2608),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1679),
            .lcout(\generator_inst1.REGSTATZ0Z_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2261),
            .ce(N__2206),
            .sr(N__2156));
    defparam \generator_inst1.REGSTAT_79_LC_2_12_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_79_LC_2_12_3 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_79_LC_2_12_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_79_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__2606),
            .in2(_gnd_net_),
            .in3(N__2018),
            .lcout(\generator_inst1.REGSTATZ0Z_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2261),
            .ce(N__2206),
            .sr(N__2156));
    defparam \generator_inst1.REGSTAT_83_LC_2_12_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_83_LC_2_12_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_83_LC_2_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_83_LC_2_12_4  (
            .in0(N__2610),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1874),
            .lcout(\generator_inst1.REGSTATZ0Z_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2261),
            .ce(N__2206),
            .sr(N__2156));
    defparam \generator_inst1.REGSTAT_2_LC_2_13_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_2_LC_2_13_0 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_2_LC_2_13_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_2_LC_2_13_0  (
            .in0(N__2586),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1904),
            .lcout(\generator_inst1.REGSTATZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2258),
            .ce(N__2204),
            .sr(N__2153));
    defparam \generator_inst1.REGSTAT_5_LC_2_13_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_5_LC_2_13_2 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_5_LC_2_13_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_5_LC_2_13_2  (
            .in0(N__2589),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1844),
            .lcout(\generator_inst1.REGSTATZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2258),
            .ce(N__2204),
            .sr(N__2153));
    defparam \generator_inst1.REGSTAT_3_LC_2_13_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_3_LC_2_13_5 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_3_LC_2_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_3_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__2587),
            .in2(_gnd_net_),
            .in3(N__1856),
            .lcout(\generator_inst1.REGSTATZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2258),
            .ce(N__2204),
            .sr(N__2153));
    defparam \generator_inst1.REGSTAT_4_LC_2_13_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_4_LC_2_13_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_4_LC_2_13_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_4_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(N__2588),
            .in2(_gnd_net_),
            .in3(N__1850),
            .lcout(\generator_inst1.REGSTATZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2258),
            .ce(N__2204),
            .sr(N__2153));
    defparam \generator_inst1.REGSTAT_25_LC_2_14_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_25_LC_2_14_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_25_LC_2_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_25_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__2578),
            .in2(_gnd_net_),
            .in3(N__1838),
            .lcout(\generator_inst1.REGSTATZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2255),
            .ce(N__2201),
            .sr(N__2150));
    defparam \generator_inst1.REGSTAT_24_LC_2_14_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_24_LC_2_14_1 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_24_LC_2_14_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_24_LC_2_14_1  (
            .in0(N__2577),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1832),
            .lcout(\generator_inst1.REGSTATZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2255),
            .ce(N__2201),
            .sr(N__2150));
    defparam \generator_inst1.REGSTAT_23_LC_2_14_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_23_LC_2_14_2 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_23_LC_2_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_23_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__2576),
            .in2(_gnd_net_),
            .in3(N__1928),
            .lcout(\generator_inst1.REGSTATZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2255),
            .ce(N__2201),
            .sr(N__2150));
    defparam \generator_inst1.REGSTAT_0_LC_2_14_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_0_LC_2_14_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_0_LC_2_14_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \generator_inst1.REGSTAT_0_LC_2_14_3  (
            .in0(N__2571),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\generator_inst1.REGSTATZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2255),
            .ce(N__2201),
            .sr(N__2150));
    defparam \generator_inst1.REGSTAT_20_LC_2_14_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_20_LC_2_14_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_20_LC_2_14_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_20_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__2573),
            .in2(_gnd_net_),
            .in3(N__1934),
            .lcout(\generator_inst1.REGSTATZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2255),
            .ce(N__2201),
            .sr(N__2150));
    defparam \generator_inst1.REGSTAT_22_LC_2_14_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_22_LC_2_14_5 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_22_LC_2_14_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_22_LC_2_14_5  (
            .in0(N__2575),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1916),
            .lcout(\generator_inst1.REGSTATZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2255),
            .ce(N__2201),
            .sr(N__2150));
    defparam \generator_inst1.REGSTAT_21_LC_2_14_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_21_LC_2_14_6 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_21_LC_2_14_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_21_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(N__2574),
            .in2(_gnd_net_),
            .in3(N__1922),
            .lcout(\generator_inst1.REGSTATZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2255),
            .ce(N__2201),
            .sr(N__2150));
    defparam \generator_inst1.REGSTAT_1_LC_2_14_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_1_LC_2_14_7 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_1_LC_2_14_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_1_LC_2_14_7  (
            .in0(N__2572),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1910),
            .lcout(\generator_inst1.REGSTATZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2255),
            .ce(N__2201),
            .sr(N__2150));
    defparam \generator_inst1.REGSTAT_30_LC_2_15_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_30_LC_2_15_0 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_30_LC_2_15_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_30_LC_2_15_0  (
            .in0(N__2569),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1886),
            .lcout(\generator_inst1.REGSTATZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2252),
            .ce(N__2198),
            .sr(N__2148));
    defparam \generator_inst1.REGSTAT_27_LC_2_15_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_27_LC_2_15_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_27_LC_2_15_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_27_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__2566),
            .in2(_gnd_net_),
            .in3(N__1988),
            .lcout(\generator_inst1.REGSTATZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2252),
            .ce(N__2198),
            .sr(N__2148));
    defparam \generator_inst1.REGSTAT_28_LC_2_15_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_28_LC_2_15_2 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_28_LC_2_15_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_28_LC_2_15_2  (
            .in0(N__2567),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1898),
            .lcout(\generator_inst1.REGSTATZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2252),
            .ce(N__2198),
            .sr(N__2148));
    defparam \generator_inst1.REGSTAT_29_LC_2_15_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_29_LC_2_15_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_29_LC_2_15_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_29_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__2568),
            .in2(_gnd_net_),
            .in3(N__1892),
            .lcout(\generator_inst1.REGSTATZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2252),
            .ce(N__2198),
            .sr(N__2148));
    defparam \generator_inst1.REGSTAT_26_LC_2_15_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_26_LC_2_15_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_26_LC_2_15_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_26_LC_2_15_4  (
            .in0(N__2565),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1994),
            .lcout(\generator_inst1.REGSTATZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2252),
            .ce(N__2198),
            .sr(N__2148));
    defparam \generator_inst1.REGSTAT_31_LC_2_15_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_31_LC_2_15_5 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_31_LC_2_15_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_31_LC_2_15_5  (
            .in0(_gnd_net_),
            .in1(N__2570),
            .in2(_gnd_net_),
            .in3(N__1982),
            .lcout(\generator_inst1.REGSTATZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2252),
            .ce(N__2198),
            .sr(N__2148));
    defparam \generator_inst1.REGSTAT_51_LC_2_16_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_51_LC_2_16_0 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_51_LC_2_16_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_51_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__2377),
            .in2(_gnd_net_),
            .in3(N__2036),
            .lcout(\generator_inst1.REGSTATZ0Z_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2250),
            .ce(N__2196),
            .sr(N__2144));
    defparam \generator_inst1.REGSTAT_47_LC_2_16_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_47_LC_2_16_1 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_47_LC_2_16_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_47_LC_2_16_1  (
            .in0(N__2373),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1952),
            .lcout(\generator_inst1.REGSTATZ0Z_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2250),
            .ce(N__2196),
            .sr(N__2144));
    defparam \generator_inst1.REGSTAT_53_LC_2_16_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_53_LC_2_16_2 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_53_LC_2_16_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_53_LC_2_16_2  (
            .in0(_gnd_net_),
            .in1(N__2379),
            .in2(_gnd_net_),
            .in3(N__1964),
            .lcout(\generator_inst1.REGSTATZ0Z_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2250),
            .ce(N__2196),
            .sr(N__2144));
    defparam \generator_inst1.REGSTAT_52_LC_2_16_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_52_LC_2_16_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_52_LC_2_16_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_52_LC_2_16_3  (
            .in0(N__2378),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1970),
            .lcout(\generator_inst1.REGSTATZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2250),
            .ce(N__2196),
            .sr(N__2144));
    defparam \generator_inst1.REGSTAT_46_LC_2_16_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_46_LC_2_16_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_46_LC_2_16_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_46_LC_2_16_4  (
            .in0(_gnd_net_),
            .in1(N__2372),
            .in2(_gnd_net_),
            .in3(N__1958),
            .lcout(\generator_inst1.REGSTATZ0Z_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2250),
            .ce(N__2196),
            .sr(N__2144));
    defparam \generator_inst1.REGSTAT_49_LC_2_16_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_49_LC_2_16_5 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_49_LC_2_16_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_49_LC_2_16_5  (
            .in0(N__2375),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1940),
            .lcout(\generator_inst1.REGSTATZ0Z_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2250),
            .ce(N__2196),
            .sr(N__2144));
    defparam \generator_inst1.REGSTAT_48_LC_2_16_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_48_LC_2_16_6 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_48_LC_2_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_48_LC_2_16_6  (
            .in0(_gnd_net_),
            .in1(N__2374),
            .in2(_gnd_net_),
            .in3(N__1946),
            .lcout(\generator_inst1.REGSTATZ0Z_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2250),
            .ce(N__2196),
            .sr(N__2144));
    defparam \generator_inst1.REGSTAT_50_LC_2_16_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_50_LC_2_16_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_50_LC_2_16_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_50_LC_2_16_7  (
            .in0(N__2376),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2042),
            .lcout(\generator_inst1.REGSTATZ0Z_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2250),
            .ce(N__2196),
            .sr(N__2144));
    defparam \generator_inst1.REGSTAT_76_LC_3_13_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_76_LC_3_13_0 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_76_LC_3_13_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_76_LC_3_13_0  (
            .in0(N__2599),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2012),
            .lcout(\generator_inst1.REGSTATZ0Z_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2262),
            .ce(N__2207),
            .sr(N__2157));
    defparam \generator_inst1.REGSTAT_77_LC_3_13_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_77_LC_3_13_1 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_77_LC_3_13_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_77_LC_3_13_1  (
            .in0(_gnd_net_),
            .in1(N__2600),
            .in2(_gnd_net_),
            .in3(N__2030),
            .lcout(\generator_inst1.REGSTATZ0Z_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2262),
            .ce(N__2207),
            .sr(N__2157));
    defparam \generator_inst1.REGSTAT_78_LC_3_13_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_78_LC_3_13_2 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_78_LC_3_13_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_78_LC_3_13_2  (
            .in0(N__2601),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2024),
            .lcout(\generator_inst1.REGSTATZ0Z_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2262),
            .ce(N__2207),
            .sr(N__2157));
    defparam \generator_inst1.REGSTAT_75_LC_3_13_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_75_LC_3_13_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_75_LC_3_13_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_75_LC_3_13_4  (
            .in0(N__2598),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2006),
            .lcout(\generator_inst1.REGSTATZ0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2262),
            .ce(N__2207),
            .sr(N__2157));
    defparam \generator_inst1.REGSTAT_74_LC_3_13_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_74_LC_3_13_7 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_74_LC_3_13_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_74_LC_3_13_7  (
            .in0(_gnd_net_),
            .in1(N__2597),
            .in2(_gnd_net_),
            .in3(N__2000),
            .lcout(\generator_inst1.REGSTATZ0Z_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2262),
            .ce(N__2207),
            .sr(N__2157));
    defparam \generator_inst1.REGSTAT_68_LC_3_14_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_68_LC_3_14_1 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_68_LC_3_14_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_68_LC_3_14_1  (
            .in0(N__2591),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2102),
            .lcout(\generator_inst1.REGSTATZ0Z_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2259),
            .ce(N__2205),
            .sr(N__2154));
    defparam \generator_inst1.REGSTAT_71_LC_3_14_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_71_LC_3_14_2 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_71_LC_3_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_71_LC_3_14_2  (
            .in0(_gnd_net_),
            .in1(N__2594),
            .in2(_gnd_net_),
            .in3(N__2096),
            .lcout(\generator_inst1.REGSTATZ0Z_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2259),
            .ce(N__2205),
            .sr(N__2154));
    defparam \generator_inst1.REGSTAT_73_LC_3_14_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_73_LC_3_14_3 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_73_LC_3_14_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_73_LC_3_14_3  (
            .in0(N__2596),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2072),
            .lcout(\generator_inst1.REGSTATZ0Z_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2259),
            .ce(N__2205),
            .sr(N__2154));
    defparam \generator_inst1.REGSTAT_67_LC_3_14_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_67_LC_3_14_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_67_LC_3_14_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_67_LC_3_14_4  (
            .in0(_gnd_net_),
            .in1(N__2590),
            .in2(_gnd_net_),
            .in3(N__2660),
            .lcout(\generator_inst1.REGSTATZ0Z_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2259),
            .ce(N__2205),
            .sr(N__2154));
    defparam \generator_inst1.REGSTAT_70_LC_3_14_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_70_LC_3_14_5 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_70_LC_3_14_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_70_LC_3_14_5  (
            .in0(N__2593),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2084),
            .lcout(\generator_inst1.REGSTATZ0Z_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2259),
            .ce(N__2205),
            .sr(N__2154));
    defparam \generator_inst1.REGSTAT_69_LC_3_14_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_69_LC_3_14_6 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_69_LC_3_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_69_LC_3_14_6  (
            .in0(_gnd_net_),
            .in1(N__2592),
            .in2(_gnd_net_),
            .in3(N__2090),
            .lcout(\generator_inst1.REGSTATZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2259),
            .ce(N__2205),
            .sr(N__2154));
    defparam \generator_inst1.REGSTAT_72_LC_3_14_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_72_LC_3_14_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_72_LC_3_14_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_72_LC_3_14_7  (
            .in0(N__2595),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2078),
            .lcout(\generator_inst1.REGSTATZ0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2259),
            .ce(N__2205),
            .sr(N__2154));
    defparam \generator_inst1.REGSTAT_64_LC_3_15_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_64_LC_3_15_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_64_LC_3_15_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_64_LC_3_15_0  (
            .in0(N__2583),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2066),
            .lcout(\generator_inst1.REGSTATZ0Z_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2256),
            .ce(N__2202),
            .sr(N__2151));
    defparam \generator_inst1.REGSTAT_60_LC_3_15_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_60_LC_3_15_1 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_60_LC_3_15_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_60_LC_3_15_1  (
            .in0(_gnd_net_),
            .in1(N__2579),
            .in2(_gnd_net_),
            .in3(N__2630),
            .lcout(\generator_inst1.REGSTATZ0Z_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2256),
            .ce(N__2202),
            .sr(N__2151));
    defparam \generator_inst1.REGSTAT_63_LC_3_15_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_63_LC_3_15_2 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_63_LC_3_15_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_63_LC_3_15_2  (
            .in0(N__2582),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2060),
            .lcout(\generator_inst1.REGSTATZ0Z_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2256),
            .ce(N__2202),
            .sr(N__2151));
    defparam \generator_inst1.REGSTAT_62_LC_3_15_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_62_LC_3_15_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_62_LC_3_15_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_62_LC_3_15_3  (
            .in0(_gnd_net_),
            .in1(N__2581),
            .in2(_gnd_net_),
            .in3(N__2048),
            .lcout(\generator_inst1.REGSTATZ0Z_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2256),
            .ce(N__2202),
            .sr(N__2151));
    defparam \generator_inst1.REGSTAT_61_LC_3_15_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_61_LC_3_15_4 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_61_LC_3_15_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_61_LC_3_15_4  (
            .in0(N__2580),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2054),
            .lcout(\generator_inst1.REGSTATZ0Z_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2256),
            .ce(N__2202),
            .sr(N__2151));
    defparam \generator_inst1.REGSTAT_66_LC_3_15_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_66_LC_3_15_5 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_66_LC_3_15_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \generator_inst1.REGSTAT_66_LC_3_15_5  (
            .in0(_gnd_net_),
            .in1(N__2585),
            .in2(_gnd_net_),
            .in3(N__2648),
            .lcout(\generator_inst1.REGSTATZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2256),
            .ce(N__2202),
            .sr(N__2151));
    defparam \generator_inst1.REGSTAT_65_LC_3_15_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_65_LC_3_15_6 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_65_LC_3_15_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_65_LC_3_15_6  (
            .in0(N__2584),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2654),
            .lcout(\generator_inst1.REGSTATZ0Z_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2256),
            .ce(N__2202),
            .sr(N__2151));
    defparam \generator_inst1.REGSTAT_57_LC_3_16_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_57_LC_3_16_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_57_LC_3_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_57_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(N__2383),
            .in2(_gnd_net_),
            .in3(N__2270),
            .lcout(\generator_inst1.REGSTATZ0Z_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2253),
            .ce(N__2199),
            .sr(N__2146));
    defparam \generator_inst1.REGSTAT_55_LC_3_16_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_55_LC_3_16_1 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_55_LC_3_16_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_55_LC_3_16_1  (
            .in0(N__2381),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2618),
            .lcout(\generator_inst1.REGSTATZ0Z_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2253),
            .ce(N__2199),
            .sr(N__2146));
    defparam \generator_inst1.REGSTAT_58_LC_3_16_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_58_LC_3_16_2 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_58_LC_3_16_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_58_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(N__2384),
            .in2(_gnd_net_),
            .in3(N__2642),
            .lcout(\generator_inst1.REGSTATZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2253),
            .ce(N__2199),
            .sr(N__2146));
    defparam \generator_inst1.REGSTAT_59_LC_3_16_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_59_LC_3_16_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_59_LC_3_16_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \generator_inst1.REGSTAT_59_LC_3_16_3  (
            .in0(N__2385),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2636),
            .lcout(\generator_inst1.REGSTATZ0Z_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2253),
            .ce(N__2199),
            .sr(N__2146));
    defparam \generator_inst1.REGSTAT_54_LC_3_16_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_54_LC_3_16_6 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_54_LC_3_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \generator_inst1.REGSTAT_54_LC_3_16_6  (
            .in0(_gnd_net_),
            .in1(N__2380),
            .in2(_gnd_net_),
            .in3(N__2624),
            .lcout(\generator_inst1.REGSTATZ0Z_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2253),
            .ce(N__2199),
            .sr(N__2146));
    defparam \generator_inst1.REGSTAT_56_LC_3_16_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_56_LC_3_16_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_56_LC_3_16_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \generator_inst1.REGSTAT_56_LC_3_16_7  (
            .in0(N__2382),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2276),
            .lcout(\generator_inst1.REGSTATZ0Z_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2253),
            .ce(N__2199),
            .sr(N__2146));
endmodule // top
