// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 12 2025 16:45:17

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    signal_out,
    RST_N,
    CLK);

    output signal_out;
    input RST_N;
    input CLK;

    wire N__1397;
    wire N__1396;
    wire N__1395;
    wire N__1388;
    wire N__1387;
    wire N__1386;
    wire N__1379;
    wire N__1378;
    wire N__1377;
    wire N__1360;
    wire N__1357;
    wire N__1354;
    wire N__1353;
    wire N__1350;
    wire N__1347;
    wire N__1342;
    wire N__1339;
    wire N__1336;
    wire N__1333;
    wire N__1332;
    wire N__1329;
    wire N__1326;
    wire N__1321;
    wire N__1318;
    wire N__1315;
    wire N__1312;
    wire N__1309;
    wire N__1308;
    wire N__1305;
    wire N__1302;
    wire N__1299;
    wire N__1294;
    wire N__1293;
    wire N__1290;
    wire N__1287;
    wire N__1284;
    wire N__1281;
    wire N__1276;
    wire N__1275;
    wire N__1272;
    wire N__1269;
    wire N__1266;
    wire N__1263;
    wire N__1258;
    wire N__1257;
    wire N__1254;
    wire N__1251;
    wire N__1248;
    wire N__1245;
    wire N__1240;
    wire N__1239;
    wire N__1236;
    wire N__1233;
    wire N__1230;
    wire N__1227;
    wire N__1222;
    wire N__1221;
    wire N__1220;
    wire N__1219;
    wire N__1218;
    wire N__1217;
    wire N__1216;
    wire N__1215;
    wire N__1214;
    wire N__1209;
    wire N__1194;
    wire N__1191;
    wire N__1188;
    wire N__1183;
    wire N__1182;
    wire N__1181;
    wire N__1178;
    wire N__1175;
    wire N__1172;
    wire N__1169;
    wire N__1166;
    wire N__1163;
    wire N__1156;
    wire N__1155;
    wire N__1154;
    wire N__1153;
    wire N__1152;
    wire N__1151;
    wire N__1138;
    wire N__1135;
    wire N__1132;
    wire N__1131;
    wire N__1130;
    wire N__1129;
    wire N__1128;
    wire N__1127;
    wire N__1114;
    wire N__1111;
    wire N__1108;
    wire N__1107;
    wire N__1104;
    wire N__1101;
    wire N__1096;
    wire N__1095;
    wire N__1094;
    wire N__1091;
    wire N__1088;
    wire N__1085;
    wire N__1078;
    wire N__1075;
    wire N__1074;
    wire N__1071;
    wire N__1068;
    wire N__1063;
    wire N__1062;
    wire N__1059;
    wire N__1056;
    wire N__1053;
    wire N__1048;
    wire N__1045;
    wire N__1042;
    wire N__1039;
    wire N__1036;
    wire N__1033;
    wire N__1030;
    wire N__1027;
    wire N__1024;
    wire N__1021;
    wire N__1018;
    wire N__1015;
    wire N__1012;
    wire N__1009;
    wire N__1006;
    wire N__1003;
    wire N__1000;
    wire N__999;
    wire N__996;
    wire N__993;
    wire N__990;
    wire N__987;
    wire N__982;
    wire N__979;
    wire N__976;
    wire N__973;
    wire N__972;
    wire N__969;
    wire N__966;
    wire N__961;
    wire N__958;
    wire N__957;
    wire N__954;
    wire N__951;
    wire N__948;
    wire N__943;
    wire N__940;
    wire N__937;
    wire N__934;
    wire N__931;
    wire N__930;
    wire N__927;
    wire N__924;
    wire N__921;
    wire N__916;
    wire N__913;
    wire N__910;
    wire N__907;
    wire N__904;
    wire N__903;
    wire N__900;
    wire N__897;
    wire N__894;
    wire N__891;
    wire N__886;
    wire N__883;
    wire N__880;
    wire N__877;
    wire N__874;
    wire N__873;
    wire N__870;
    wire N__867;
    wire N__862;
    wire N__859;
    wire N__856;
    wire N__855;
    wire N__852;
    wire N__849;
    wire N__844;
    wire N__841;
    wire N__840;
    wire N__837;
    wire N__834;
    wire N__829;
    wire N__826;
    wire N__825;
    wire N__822;
    wire N__819;
    wire N__814;
    wire N__811;
    wire N__810;
    wire N__807;
    wire N__804;
    wire N__801;
    wire N__798;
    wire N__793;
    wire N__790;
    wire N__787;
    wire N__784;
    wire N__781;
    wire N__780;
    wire N__777;
    wire N__774;
    wire N__769;
    wire N__766;
    wire N__763;
    wire N__762;
    wire N__759;
    wire N__756;
    wire N__751;
    wire N__748;
    wire N__745;
    wire N__742;
    wire N__739;
    wire N__738;
    wire N__737;
    wire N__736;
    wire N__735;
    wire N__734;
    wire N__733;
    wire N__732;
    wire N__731;
    wire N__716;
    wire N__711;
    wire N__706;
    wire N__705;
    wire N__704;
    wire N__703;
    wire N__702;
    wire N__701;
    wire N__698;
    wire N__697;
    wire N__694;
    wire N__693;
    wire N__692;
    wire N__689;
    wire N__686;
    wire N__683;
    wire N__680;
    wire N__677;
    wire N__672;
    wire N__659;
    wire N__652;
    wire N__651;
    wire N__646;
    wire N__643;
    wire N__640;
    wire N__637;
    wire N__634;
    wire N__631;
    wire N__628;
    wire N__625;
    wire N__622;
    wire N__619;
    wire N__616;
    wire N__613;
    wire N__610;
    wire N__607;
    wire N__604;
    wire N__601;
    wire N__598;
    wire N__595;
    wire N__592;
    wire N__589;
    wire N__586;
    wire N__583;
    wire CLK_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \generator_inst1.signal_out5_11 ;
    wire \generator_inst1.signal_out5_13_cascade_ ;
    wire \generator_inst1.signal_out5_14 ;
    wire \generator_inst1.signal_out5_15 ;
    wire \generator_inst1.signal_out5_20 ;
    wire generated_signal;
    wire signal_out_c;
    wire bfn_11_17_0_;
    wire \generator_inst1.un3_counter_1_cry_1 ;
    wire \generator_inst1.un3_counter_1_cry_2 ;
    wire \generator_inst1.un3_counter_1_cry_3 ;
    wire \generator_inst1.counterZ0Z_5 ;
    wire \generator_inst1.un3_counter_1_cry_4 ;
    wire \generator_inst1.counterZ0Z_6 ;
    wire \generator_inst1.un3_counter_1_cry_5 ;
    wire \generator_inst1.counterZ0Z_7 ;
    wire \generator_inst1.un3_counter_1_cry_6 ;
    wire \generator_inst1.counterZ0Z_8 ;
    wire \generator_inst1.un3_counter_1_cry_7 ;
    wire \generator_inst1.un3_counter_1_cry_8 ;
    wire \generator_inst1.counterZ0Z_9 ;
    wire \generator_inst1.counter_RNO_0Z0Z_9 ;
    wire bfn_11_18_0_;
    wire \generator_inst1.counterZ0Z_10 ;
    wire \generator_inst1.un3_counter_1_cry_9 ;
    wire \generator_inst1.un3_counter_1_cry_10 ;
    wire \generator_inst1.counterZ0Z_12 ;
    wire \generator_inst1.counter_RNO_0Z0Z_12 ;
    wire \generator_inst1.un3_counter_1_cry_11 ;
    wire \generator_inst1.counterZ0Z_13 ;
    wire \generator_inst1.un3_counter_1_cry_12 ;
    wire \generator_inst1.un3_counter_1_cry_13 ;
    wire \generator_inst1.un3_counter_1_cry_14 ;
    wire \generator_inst1.counterZ0Z_16 ;
    wire \generator_inst1.un3_counter_1_cry_15 ;
    wire \generator_inst1.un3_counter_1_cry_16 ;
    wire \generator_inst1.counterZ0Z_17 ;
    wire \generator_inst1.counter_RNO_0Z0Z_17 ;
    wire bfn_11_19_0_;
    wire \generator_inst1.un3_counter_1_cry_17 ;
    wire \generator_inst1.counterZ0Z_19 ;
    wire \generator_inst1.counter_RNO_0Z0Z_19 ;
    wire \generator_inst1.un3_counter_1_cry_18 ;
    wire \generator_inst1.counterZ0Z_20 ;
    wire \generator_inst1.counter_RNO_0Z0Z_20 ;
    wire \generator_inst1.un3_counter_1_cry_19 ;
    wire \generator_inst1.counterZ0Z_21 ;
    wire \generator_inst1.counter_RNO_0Z0Z_21 ;
    wire \generator_inst1.un3_counter_1_cry_20 ;
    wire \generator_inst1.counterZ0Z_22 ;
    wire \generator_inst1.counter_RNO_0Z0Z_22 ;
    wire \generator_inst1.un3_counter_1_cry_21 ;
    wire \generator_inst1.un3_counter_1_cry_22 ;
    wire \generator_inst1.counterZ0Z_23 ;
    wire \generator_inst1.counterZ0Z_11 ;
    wire \generator_inst1.counterZ0Z_3 ;
    wire \generator_inst1.counterZ0Z_18 ;
    wire \generator_inst1.counterZ0Z_2 ;
    wire \generator_inst1.signal_out5_16 ;
    wire \generator_inst1.counterZ0Z_0 ;
    wire CLK_c_g;
    wire RST_N_c_i_g;
    wire \generator_inst1.counterZ0Z_4 ;
    wire \generator_inst1.counterZ0Z_1 ;
    wire \generator_inst1.counterZ0Z_14 ;
    wire \generator_inst1.counterZ0Z_15 ;
    wire \generator_inst1.signal_out5_12 ;
    wire RST_N_c;
    wire RST_N_c_i;
    wire _gnd_net_;

    IO_PAD RST_N_ibuf_iopad (
            .OE(N__1397),
            .DIN(N__1396),
            .DOUT(N__1395),
            .PACKAGEPIN(RST_N));
    defparam RST_N_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RST_N_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RST_N_ibuf_preio (
            .PADOEN(N__1397),
            .PADOUT(N__1396),
            .PADIN(N__1395),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RST_N_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD signal_out_obuf_iopad (
            .OE(N__1388),
            .DIN(N__1387),
            .DOUT(N__1386),
            .PACKAGEPIN(signal_out));
    defparam signal_out_obuf_preio.NEG_TRIGGER=1'b0;
    defparam signal_out_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO signal_out_obuf_preio (
            .PADOEN(N__1388),
            .PADOUT(N__1387),
            .PADIN(N__1386),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__643),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__1379),
            .DIN(N__1378),
            .DOUT(N__1377),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__1379),
            .PADOUT(N__1378),
            .PADIN(N__1377),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__312 (
            .O(N__1360),
            .I(N__1357));
    InMux I__311 (
            .O(N__1357),
            .I(N__1354));
    LocalMux I__310 (
            .O(N__1354),
            .I(N__1350));
    InMux I__309 (
            .O(N__1353),
            .I(N__1347));
    Odrv12 I__308 (
            .O(N__1350),
            .I(\generator_inst1.counterZ0Z_21 ));
    LocalMux I__307 (
            .O(N__1347),
            .I(\generator_inst1.counterZ0Z_21 ));
    InMux I__306 (
            .O(N__1342),
            .I(N__1339));
    LocalMux I__305 (
            .O(N__1339),
            .I(\generator_inst1.counter_RNO_0Z0Z_21 ));
    InMux I__304 (
            .O(N__1336),
            .I(\generator_inst1.un3_counter_1_cry_20 ));
    InMux I__303 (
            .O(N__1333),
            .I(N__1329));
    InMux I__302 (
            .O(N__1332),
            .I(N__1326));
    LocalMux I__301 (
            .O(N__1329),
            .I(\generator_inst1.counterZ0Z_22 ));
    LocalMux I__300 (
            .O(N__1326),
            .I(\generator_inst1.counterZ0Z_22 ));
    InMux I__299 (
            .O(N__1321),
            .I(N__1318));
    LocalMux I__298 (
            .O(N__1318),
            .I(\generator_inst1.counter_RNO_0Z0Z_22 ));
    InMux I__297 (
            .O(N__1315),
            .I(\generator_inst1.un3_counter_1_cry_21 ));
    InMux I__296 (
            .O(N__1312),
            .I(\generator_inst1.un3_counter_1_cry_22 ));
    CascadeMux I__295 (
            .O(N__1309),
            .I(N__1305));
    InMux I__294 (
            .O(N__1308),
            .I(N__1302));
    InMux I__293 (
            .O(N__1305),
            .I(N__1299));
    LocalMux I__292 (
            .O(N__1302),
            .I(\generator_inst1.counterZ0Z_23 ));
    LocalMux I__291 (
            .O(N__1299),
            .I(\generator_inst1.counterZ0Z_23 ));
    InMux I__290 (
            .O(N__1294),
            .I(N__1290));
    CascadeMux I__289 (
            .O(N__1293),
            .I(N__1287));
    LocalMux I__288 (
            .O(N__1290),
            .I(N__1284));
    InMux I__287 (
            .O(N__1287),
            .I(N__1281));
    Odrv4 I__286 (
            .O(N__1284),
            .I(\generator_inst1.counterZ0Z_11 ));
    LocalMux I__285 (
            .O(N__1281),
            .I(\generator_inst1.counterZ0Z_11 ));
    InMux I__284 (
            .O(N__1276),
            .I(N__1272));
    CascadeMux I__283 (
            .O(N__1275),
            .I(N__1269));
    LocalMux I__282 (
            .O(N__1272),
            .I(N__1266));
    InMux I__281 (
            .O(N__1269),
            .I(N__1263));
    Odrv4 I__280 (
            .O(N__1266),
            .I(\generator_inst1.counterZ0Z_3 ));
    LocalMux I__279 (
            .O(N__1263),
            .I(\generator_inst1.counterZ0Z_3 ));
    CascadeMux I__278 (
            .O(N__1258),
            .I(N__1254));
    CascadeMux I__277 (
            .O(N__1257),
            .I(N__1251));
    InMux I__276 (
            .O(N__1254),
            .I(N__1248));
    InMux I__275 (
            .O(N__1251),
            .I(N__1245));
    LocalMux I__274 (
            .O(N__1248),
            .I(\generator_inst1.counterZ0Z_18 ));
    LocalMux I__273 (
            .O(N__1245),
            .I(\generator_inst1.counterZ0Z_18 ));
    InMux I__272 (
            .O(N__1240),
            .I(N__1236));
    CascadeMux I__271 (
            .O(N__1239),
            .I(N__1233));
    LocalMux I__270 (
            .O(N__1236),
            .I(N__1230));
    InMux I__269 (
            .O(N__1233),
            .I(N__1227));
    Odrv12 I__268 (
            .O(N__1230),
            .I(\generator_inst1.counterZ0Z_2 ));
    LocalMux I__267 (
            .O(N__1227),
            .I(\generator_inst1.counterZ0Z_2 ));
    InMux I__266 (
            .O(N__1222),
            .I(N__1209));
    InMux I__265 (
            .O(N__1221),
            .I(N__1209));
    InMux I__264 (
            .O(N__1220),
            .I(N__1194));
    InMux I__263 (
            .O(N__1219),
            .I(N__1194));
    InMux I__262 (
            .O(N__1218),
            .I(N__1194));
    InMux I__261 (
            .O(N__1217),
            .I(N__1194));
    InMux I__260 (
            .O(N__1216),
            .I(N__1194));
    InMux I__259 (
            .O(N__1215),
            .I(N__1194));
    InMux I__258 (
            .O(N__1214),
            .I(N__1194));
    LocalMux I__257 (
            .O(N__1209),
            .I(N__1191));
    LocalMux I__256 (
            .O(N__1194),
            .I(N__1188));
    Odrv4 I__255 (
            .O(N__1191),
            .I(\generator_inst1.signal_out5_16 ));
    Odrv4 I__254 (
            .O(N__1188),
            .I(\generator_inst1.signal_out5_16 ));
    CascadeMux I__253 (
            .O(N__1183),
            .I(N__1178));
    InMux I__252 (
            .O(N__1182),
            .I(N__1175));
    CascadeMux I__251 (
            .O(N__1181),
            .I(N__1172));
    InMux I__250 (
            .O(N__1178),
            .I(N__1169));
    LocalMux I__249 (
            .O(N__1175),
            .I(N__1166));
    InMux I__248 (
            .O(N__1172),
            .I(N__1163));
    LocalMux I__247 (
            .O(N__1169),
            .I(\generator_inst1.counterZ0Z_0 ));
    Odrv4 I__246 (
            .O(N__1166),
            .I(\generator_inst1.counterZ0Z_0 ));
    LocalMux I__245 (
            .O(N__1163),
            .I(\generator_inst1.counterZ0Z_0 ));
    ClkMux I__244 (
            .O(N__1156),
            .I(N__1138));
    ClkMux I__243 (
            .O(N__1155),
            .I(N__1138));
    ClkMux I__242 (
            .O(N__1154),
            .I(N__1138));
    ClkMux I__241 (
            .O(N__1153),
            .I(N__1138));
    ClkMux I__240 (
            .O(N__1152),
            .I(N__1138));
    ClkMux I__239 (
            .O(N__1151),
            .I(N__1138));
    GlobalMux I__238 (
            .O(N__1138),
            .I(N__1135));
    gio2CtrlBuf I__237 (
            .O(N__1135),
            .I(CLK_c_g));
    SRMux I__236 (
            .O(N__1132),
            .I(N__1114));
    SRMux I__235 (
            .O(N__1131),
            .I(N__1114));
    SRMux I__234 (
            .O(N__1130),
            .I(N__1114));
    SRMux I__233 (
            .O(N__1129),
            .I(N__1114));
    SRMux I__232 (
            .O(N__1128),
            .I(N__1114));
    SRMux I__231 (
            .O(N__1127),
            .I(N__1114));
    GlobalMux I__230 (
            .O(N__1114),
            .I(N__1111));
    gio2CtrlBuf I__229 (
            .O(N__1111),
            .I(RST_N_c_i_g));
    InMux I__228 (
            .O(N__1108),
            .I(N__1104));
    InMux I__227 (
            .O(N__1107),
            .I(N__1101));
    LocalMux I__226 (
            .O(N__1104),
            .I(\generator_inst1.counterZ0Z_4 ));
    LocalMux I__225 (
            .O(N__1101),
            .I(\generator_inst1.counterZ0Z_4 ));
    InMux I__224 (
            .O(N__1096),
            .I(N__1091));
    InMux I__223 (
            .O(N__1095),
            .I(N__1088));
    InMux I__222 (
            .O(N__1094),
            .I(N__1085));
    LocalMux I__221 (
            .O(N__1091),
            .I(\generator_inst1.counterZ0Z_1 ));
    LocalMux I__220 (
            .O(N__1088),
            .I(\generator_inst1.counterZ0Z_1 ));
    LocalMux I__219 (
            .O(N__1085),
            .I(\generator_inst1.counterZ0Z_1 ));
    CascadeMux I__218 (
            .O(N__1078),
            .I(N__1075));
    InMux I__217 (
            .O(N__1075),
            .I(N__1071));
    InMux I__216 (
            .O(N__1074),
            .I(N__1068));
    LocalMux I__215 (
            .O(N__1071),
            .I(\generator_inst1.counterZ0Z_14 ));
    LocalMux I__214 (
            .O(N__1068),
            .I(\generator_inst1.counterZ0Z_14 ));
    CascadeMux I__213 (
            .O(N__1063),
            .I(N__1059));
    InMux I__212 (
            .O(N__1062),
            .I(N__1056));
    InMux I__211 (
            .O(N__1059),
            .I(N__1053));
    LocalMux I__210 (
            .O(N__1056),
            .I(\generator_inst1.counterZ0Z_15 ));
    LocalMux I__209 (
            .O(N__1053),
            .I(\generator_inst1.counterZ0Z_15 ));
    InMux I__208 (
            .O(N__1048),
            .I(N__1045));
    LocalMux I__207 (
            .O(N__1045),
            .I(N__1042));
    Odrv12 I__206 (
            .O(N__1042),
            .I(\generator_inst1.signal_out5_12 ));
    InMux I__205 (
            .O(N__1039),
            .I(N__1036));
    LocalMux I__204 (
            .O(N__1036),
            .I(N__1033));
    Span12Mux_v I__203 (
            .O(N__1033),
            .I(N__1030));
    Odrv12 I__202 (
            .O(N__1030),
            .I(RST_N_c));
    IoInMux I__201 (
            .O(N__1027),
            .I(N__1024));
    LocalMux I__200 (
            .O(N__1024),
            .I(N__1021));
    Span4Mux_s1_h I__199 (
            .O(N__1021),
            .I(N__1018));
    Span4Mux_h I__198 (
            .O(N__1018),
            .I(N__1015));
    Sp12to4 I__197 (
            .O(N__1015),
            .I(N__1012));
    Span12Mux_v I__196 (
            .O(N__1012),
            .I(N__1009));
    Span12Mux_h I__195 (
            .O(N__1009),
            .I(N__1006));
    Span12Mux_h I__194 (
            .O(N__1006),
            .I(N__1003));
    Odrv12 I__193 (
            .O(N__1003),
            .I(RST_N_c_i));
    CascadeMux I__192 (
            .O(N__1000),
            .I(N__996));
    CascadeMux I__191 (
            .O(N__999),
            .I(N__993));
    InMux I__190 (
            .O(N__996),
            .I(N__990));
    InMux I__189 (
            .O(N__993),
            .I(N__987));
    LocalMux I__188 (
            .O(N__990),
            .I(\generator_inst1.counterZ0Z_13 ));
    LocalMux I__187 (
            .O(N__987),
            .I(\generator_inst1.counterZ0Z_13 ));
    InMux I__186 (
            .O(N__982),
            .I(\generator_inst1.un3_counter_1_cry_12 ));
    InMux I__185 (
            .O(N__979),
            .I(\generator_inst1.un3_counter_1_cry_13 ));
    InMux I__184 (
            .O(N__976),
            .I(\generator_inst1.un3_counter_1_cry_14 ));
    InMux I__183 (
            .O(N__973),
            .I(N__969));
    InMux I__182 (
            .O(N__972),
            .I(N__966));
    LocalMux I__181 (
            .O(N__969),
            .I(\generator_inst1.counterZ0Z_16 ));
    LocalMux I__180 (
            .O(N__966),
            .I(\generator_inst1.counterZ0Z_16 ));
    InMux I__179 (
            .O(N__961),
            .I(\generator_inst1.un3_counter_1_cry_15 ));
    InMux I__178 (
            .O(N__958),
            .I(N__954));
    InMux I__177 (
            .O(N__957),
            .I(N__951));
    LocalMux I__176 (
            .O(N__954),
            .I(N__948));
    LocalMux I__175 (
            .O(N__951),
            .I(\generator_inst1.counterZ0Z_17 ));
    Odrv4 I__174 (
            .O(N__948),
            .I(\generator_inst1.counterZ0Z_17 ));
    InMux I__173 (
            .O(N__943),
            .I(N__940));
    LocalMux I__172 (
            .O(N__940),
            .I(\generator_inst1.counter_RNO_0Z0Z_17 ));
    InMux I__171 (
            .O(N__937),
            .I(bfn_11_19_0_));
    InMux I__170 (
            .O(N__934),
            .I(\generator_inst1.un3_counter_1_cry_17 ));
    CascadeMux I__169 (
            .O(N__931),
            .I(N__927));
    InMux I__168 (
            .O(N__930),
            .I(N__924));
    InMux I__167 (
            .O(N__927),
            .I(N__921));
    LocalMux I__166 (
            .O(N__924),
            .I(\generator_inst1.counterZ0Z_19 ));
    LocalMux I__165 (
            .O(N__921),
            .I(\generator_inst1.counterZ0Z_19 ));
    CascadeMux I__164 (
            .O(N__916),
            .I(N__913));
    InMux I__163 (
            .O(N__913),
            .I(N__910));
    LocalMux I__162 (
            .O(N__910),
            .I(\generator_inst1.counter_RNO_0Z0Z_19 ));
    InMux I__161 (
            .O(N__907),
            .I(\generator_inst1.un3_counter_1_cry_18 ));
    CascadeMux I__160 (
            .O(N__904),
            .I(N__900));
    CascadeMux I__159 (
            .O(N__903),
            .I(N__897));
    InMux I__158 (
            .O(N__900),
            .I(N__894));
    InMux I__157 (
            .O(N__897),
            .I(N__891));
    LocalMux I__156 (
            .O(N__894),
            .I(\generator_inst1.counterZ0Z_20 ));
    LocalMux I__155 (
            .O(N__891),
            .I(\generator_inst1.counterZ0Z_20 ));
    InMux I__154 (
            .O(N__886),
            .I(N__883));
    LocalMux I__153 (
            .O(N__883),
            .I(\generator_inst1.counter_RNO_0Z0Z_20 ));
    InMux I__152 (
            .O(N__880),
            .I(\generator_inst1.un3_counter_1_cry_19 ));
    InMux I__151 (
            .O(N__877),
            .I(\generator_inst1.un3_counter_1_cry_3 ));
    InMux I__150 (
            .O(N__874),
            .I(N__870));
    InMux I__149 (
            .O(N__873),
            .I(N__867));
    LocalMux I__148 (
            .O(N__870),
            .I(\generator_inst1.counterZ0Z_5 ));
    LocalMux I__147 (
            .O(N__867),
            .I(\generator_inst1.counterZ0Z_5 ));
    InMux I__146 (
            .O(N__862),
            .I(\generator_inst1.un3_counter_1_cry_4 ));
    InMux I__145 (
            .O(N__859),
            .I(N__856));
    LocalMux I__144 (
            .O(N__856),
            .I(N__852));
    InMux I__143 (
            .O(N__855),
            .I(N__849));
    Odrv4 I__142 (
            .O(N__852),
            .I(\generator_inst1.counterZ0Z_6 ));
    LocalMux I__141 (
            .O(N__849),
            .I(\generator_inst1.counterZ0Z_6 ));
    InMux I__140 (
            .O(N__844),
            .I(\generator_inst1.un3_counter_1_cry_5 ));
    InMux I__139 (
            .O(N__841),
            .I(N__837));
    InMux I__138 (
            .O(N__840),
            .I(N__834));
    LocalMux I__137 (
            .O(N__837),
            .I(\generator_inst1.counterZ0Z_7 ));
    LocalMux I__136 (
            .O(N__834),
            .I(\generator_inst1.counterZ0Z_7 ));
    InMux I__135 (
            .O(N__829),
            .I(\generator_inst1.un3_counter_1_cry_6 ));
    InMux I__134 (
            .O(N__826),
            .I(N__822));
    InMux I__133 (
            .O(N__825),
            .I(N__819));
    LocalMux I__132 (
            .O(N__822),
            .I(\generator_inst1.counterZ0Z_8 ));
    LocalMux I__131 (
            .O(N__819),
            .I(\generator_inst1.counterZ0Z_8 ));
    InMux I__130 (
            .O(N__814),
            .I(\generator_inst1.un3_counter_1_cry_7 ));
    InMux I__129 (
            .O(N__811),
            .I(N__807));
    CascadeMux I__128 (
            .O(N__810),
            .I(N__804));
    LocalMux I__127 (
            .O(N__807),
            .I(N__801));
    InMux I__126 (
            .O(N__804),
            .I(N__798));
    Odrv4 I__125 (
            .O(N__801),
            .I(\generator_inst1.counterZ0Z_9 ));
    LocalMux I__124 (
            .O(N__798),
            .I(\generator_inst1.counterZ0Z_9 ));
    InMux I__123 (
            .O(N__793),
            .I(N__790));
    LocalMux I__122 (
            .O(N__790),
            .I(\generator_inst1.counter_RNO_0Z0Z_9 ));
    InMux I__121 (
            .O(N__787),
            .I(bfn_11_18_0_));
    InMux I__120 (
            .O(N__784),
            .I(N__781));
    LocalMux I__119 (
            .O(N__781),
            .I(N__777));
    InMux I__118 (
            .O(N__780),
            .I(N__774));
    Odrv4 I__117 (
            .O(N__777),
            .I(\generator_inst1.counterZ0Z_10 ));
    LocalMux I__116 (
            .O(N__774),
            .I(\generator_inst1.counterZ0Z_10 ));
    InMux I__115 (
            .O(N__769),
            .I(\generator_inst1.un3_counter_1_cry_9 ));
    InMux I__114 (
            .O(N__766),
            .I(\generator_inst1.un3_counter_1_cry_10 ));
    InMux I__113 (
            .O(N__763),
            .I(N__759));
    InMux I__112 (
            .O(N__762),
            .I(N__756));
    LocalMux I__111 (
            .O(N__759),
            .I(\generator_inst1.counterZ0Z_12 ));
    LocalMux I__110 (
            .O(N__756),
            .I(\generator_inst1.counterZ0Z_12 ));
    CascadeMux I__109 (
            .O(N__751),
            .I(N__748));
    InMux I__108 (
            .O(N__748),
            .I(N__745));
    LocalMux I__107 (
            .O(N__745),
            .I(\generator_inst1.counter_RNO_0Z0Z_12 ));
    InMux I__106 (
            .O(N__742),
            .I(\generator_inst1.un3_counter_1_cry_11 ));
    InMux I__105 (
            .O(N__739),
            .I(N__716));
    InMux I__104 (
            .O(N__738),
            .I(N__716));
    InMux I__103 (
            .O(N__737),
            .I(N__716));
    InMux I__102 (
            .O(N__736),
            .I(N__716));
    InMux I__101 (
            .O(N__735),
            .I(N__716));
    InMux I__100 (
            .O(N__734),
            .I(N__716));
    InMux I__99 (
            .O(N__733),
            .I(N__716));
    InMux I__98 (
            .O(N__732),
            .I(N__711));
    InMux I__97 (
            .O(N__731),
            .I(N__711));
    LocalMux I__96 (
            .O(N__716),
            .I(\generator_inst1.signal_out5_15 ));
    LocalMux I__95 (
            .O(N__711),
            .I(\generator_inst1.signal_out5_15 ));
    CascadeMux I__94 (
            .O(N__706),
            .I(N__698));
    CascadeMux I__93 (
            .O(N__705),
            .I(N__694));
    CascadeMux I__92 (
            .O(N__704),
            .I(N__689));
    CascadeMux I__91 (
            .O(N__703),
            .I(N__686));
    CascadeMux I__90 (
            .O(N__702),
            .I(N__683));
    CascadeMux I__89 (
            .O(N__701),
            .I(N__680));
    InMux I__88 (
            .O(N__698),
            .I(N__677));
    InMux I__87 (
            .O(N__697),
            .I(N__672));
    InMux I__86 (
            .O(N__694),
            .I(N__672));
    InMux I__85 (
            .O(N__693),
            .I(N__659));
    InMux I__84 (
            .O(N__692),
            .I(N__659));
    InMux I__83 (
            .O(N__689),
            .I(N__659));
    InMux I__82 (
            .O(N__686),
            .I(N__659));
    InMux I__81 (
            .O(N__683),
            .I(N__659));
    InMux I__80 (
            .O(N__680),
            .I(N__659));
    LocalMux I__79 (
            .O(N__677),
            .I(\generator_inst1.signal_out5_20 ));
    LocalMux I__78 (
            .O(N__672),
            .I(\generator_inst1.signal_out5_20 ));
    LocalMux I__77 (
            .O(N__659),
            .I(\generator_inst1.signal_out5_20 ));
    InMux I__76 (
            .O(N__652),
            .I(N__646));
    InMux I__75 (
            .O(N__651),
            .I(N__646));
    LocalMux I__74 (
            .O(N__646),
            .I(generated_signal));
    IoInMux I__73 (
            .O(N__643),
            .I(N__640));
    LocalMux I__72 (
            .O(N__640),
            .I(N__637));
    IoSpan4Mux I__71 (
            .O(N__637),
            .I(N__634));
    Span4Mux_s2_v I__70 (
            .O(N__634),
            .I(N__631));
    Sp12to4 I__69 (
            .O(N__631),
            .I(N__628));
    Span12Mux_v I__68 (
            .O(N__628),
            .I(N__625));
    Span12Mux_h I__67 (
            .O(N__625),
            .I(N__622));
    Odrv12 I__66 (
            .O(N__622),
            .I(signal_out_c));
    InMux I__65 (
            .O(N__619),
            .I(\generator_inst1.un3_counter_1_cry_1 ));
    InMux I__64 (
            .O(N__616),
            .I(\generator_inst1.un3_counter_1_cry_2 ));
    InMux I__63 (
            .O(N__613),
            .I(N__610));
    LocalMux I__62 (
            .O(N__610),
            .I(\generator_inst1.signal_out5_11 ));
    CascadeMux I__61 (
            .O(N__607),
            .I(\generator_inst1.signal_out5_13_cascade_ ));
    InMux I__60 (
            .O(N__604),
            .I(N__601));
    LocalMux I__59 (
            .O(N__601),
            .I(\generator_inst1.signal_out5_14 ));
    IoInMux I__58 (
            .O(N__598),
            .I(N__595));
    LocalMux I__57 (
            .O(N__595),
            .I(N__592));
    IoSpan4Mux I__56 (
            .O(N__592),
            .I(N__589));
    IoSpan4Mux I__55 (
            .O(N__589),
            .I(N__586));
    IoSpan4Mux I__54 (
            .O(N__586),
            .I(N__583));
    Odrv4 I__53 (
            .O(N__583),
            .I(CLK_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\generator_inst1.un3_counter_1_cry_8 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(\generator_inst1.un3_counter_1_cry_16 ),
            .carryinitout(bfn_11_19_0_));
    ICE_GB CLK_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__598),
            .GLOBALBUFFEROUTPUT(CLK_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB RST_N_ibuf_RNIBJGC_0 (
            .USERSIGNALTOGLOBALBUFFER(N__1027),
            .GLOBALBUFFEROUTPUT(RST_N_c_i_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \generator_inst1.counter_0_LC_10_17_3 .C_ON=1'b0;
    defparam \generator_inst1.counter_0_LC_10_17_3 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_0_LC_10_17_3 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \generator_inst1.counter_0_LC_10_17_3  (
            .in0(N__1221),
            .in1(N__731),
            .in2(N__1183),
            .in3(N__697),
            .lcout(\generator_inst1.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1151),
            .ce(),
            .sr(N__1127));
    defparam \generator_inst1.counter_9_LC_10_17_4 .C_ON=1'b0;
    defparam \generator_inst1.counter_9_LC_10_17_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_9_LC_10_17_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \generator_inst1.counter_9_LC_10_17_4  (
            .in0(N__732),
            .in1(N__1222),
            .in2(N__705),
            .in3(N__793),
            .lcout(\generator_inst1.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1151),
            .ce(),
            .sr(N__1127));
    defparam \generator_inst1.counter_RNI30RL1_12_LC_10_18_0 .C_ON=1'b0;
    defparam \generator_inst1.counter_RNI30RL1_12_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.counter_RNI30RL1_12_LC_10_18_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \generator_inst1.counter_RNI30RL1_12_LC_10_18_0  (
            .in0(N__958),
            .in1(N__763),
            .in2(N__904),
            .in3(N__930),
            .lcout(\generator_inst1.signal_out5_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.counter_RNIIF331_23_LC_10_18_1 .C_ON=1'b0;
    defparam \generator_inst1.counter_RNIIF331_23_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.counter_RNIIF331_23_LC_10_18_1 .LUT_INIT=16'b0000000100000001;
    LogicCell40 \generator_inst1.counter_RNIIF331_23_LC_10_18_1  (
            .in0(N__973),
            .in1(N__874),
            .in2(N__1309),
            .in3(_gnd_net_),
            .lcout(\generator_inst1.signal_out5_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.counter_RNIM0V51_6_LC_10_18_4 .C_ON=1'b0;
    defparam \generator_inst1.counter_RNIM0V51_6_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.counter_RNIM0V51_6_LC_10_18_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \generator_inst1.counter_RNIM0V51_6_LC_10_18_4  (
            .in0(N__811),
            .in1(N__841),
            .in2(N__1000),
            .in3(N__859),
            .lcout(\generator_inst1.signal_out5_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.counter_RNICPIG1_8_LC_10_18_5 .C_ON=1'b0;
    defparam \generator_inst1.counter_RNICPIG1_8_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.counter_RNICPIG1_8_LC_10_18_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \generator_inst1.counter_RNICPIG1_8_LC_10_18_5  (
            .in0(N__784),
            .in1(N__826),
            .in2(N__1360),
            .in3(N__1332),
            .lcout(),
            .ltout(\generator_inst1.signal_out5_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.counter_RNITVOK5_1_LC_10_18_6 .C_ON=1'b0;
    defparam \generator_inst1.counter_RNITVOK5_1_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.counter_RNITVOK5_1_LC_10_18_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \generator_inst1.counter_RNITVOK5_1_LC_10_18_6  (
            .in0(N__613),
            .in1(N__1048),
            .in2(N__607),
            .in3(N__604),
            .lcout(\generator_inst1.signal_out5_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.signal_out_LC_10_19_0 .C_ON=1'b0;
    defparam \generator_inst1.signal_out_LC_10_19_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.signal_out_LC_10_19_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \generator_inst1.signal_out_LC_10_19_0  (
            .in0(N__739),
            .in1(N__651),
            .in2(N__704),
            .in3(N__1220),
            .lcout(generated_signal),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1154),
            .ce(),
            .sr(N__1129));
    defparam \generator_inst1.counter_21_LC_10_19_1 .C_ON=1'b0;
    defparam \generator_inst1.counter_21_LC_10_19_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_21_LC_10_19_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \generator_inst1.counter_21_LC_10_19_1  (
            .in0(N__1218),
            .in1(N__737),
            .in2(N__706),
            .in3(N__1342),
            .lcout(\generator_inst1.counterZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1154),
            .ce(),
            .sr(N__1129));
    defparam \generator_inst1.counter_22_LC_10_19_2 .C_ON=1'b0;
    defparam \generator_inst1.counter_22_LC_10_19_2 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_22_LC_10_19_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \generator_inst1.counter_22_LC_10_19_2  (
            .in0(N__738),
            .in1(N__1219),
            .in2(N__703),
            .in3(N__1321),
            .lcout(\generator_inst1.counterZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1154),
            .ce(),
            .sr(N__1129));
    defparam \generator_inst1.counter_12_LC_10_19_3 .C_ON=1'b0;
    defparam \generator_inst1.counter_12_LC_10_19_3 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_12_LC_10_19_3 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \generator_inst1.counter_12_LC_10_19_3  (
            .in0(N__1214),
            .in1(N__733),
            .in2(N__751),
            .in3(N__692),
            .lcout(\generator_inst1.counterZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1154),
            .ce(),
            .sr(N__1129));
    defparam \generator_inst1.counter_17_LC_10_19_4 .C_ON=1'b0;
    defparam \generator_inst1.counter_17_LC_10_19_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_17_LC_10_19_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \generator_inst1.counter_17_LC_10_19_4  (
            .in0(N__734),
            .in1(N__1215),
            .in2(N__701),
            .in3(N__943),
            .lcout(\generator_inst1.counterZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1154),
            .ce(),
            .sr(N__1129));
    defparam \generator_inst1.counter_19_LC_10_19_5 .C_ON=1'b0;
    defparam \generator_inst1.counter_19_LC_10_19_5 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_19_LC_10_19_5 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \generator_inst1.counter_19_LC_10_19_5  (
            .in0(N__1216),
            .in1(N__735),
            .in2(N__916),
            .in3(N__693),
            .lcout(\generator_inst1.counterZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1154),
            .ce(),
            .sr(N__1129));
    defparam \generator_inst1.counter_20_LC_10_19_6 .C_ON=1'b0;
    defparam \generator_inst1.counter_20_LC_10_19_6 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_20_LC_10_19_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \generator_inst1.counter_20_LC_10_19_6  (
            .in0(N__736),
            .in1(N__1217),
            .in2(N__702),
            .in3(N__886),
            .lcout(\generator_inst1.counterZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1154),
            .ce(),
            .sr(N__1129));
    defparam \receptor_inst1.signal_out_LC_10_19_7 .C_ON=1'b0;
    defparam \receptor_inst1.signal_out_LC_10_19_7 .SEQ_MODE=4'b1010;
    defparam \receptor_inst1.signal_out_LC_10_19_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \receptor_inst1.signal_out_LC_10_19_7  (
            .in0(N__652),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(signal_out_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1154),
            .ce(),
            .sr(N__1129));
    defparam \generator_inst1.un3_counter_1_cry_1_c_LC_11_17_0 .C_ON=1'b1;
    defparam \generator_inst1.un3_counter_1_cry_1_c_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.un3_counter_1_cry_1_c_LC_11_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \generator_inst1.un3_counter_1_cry_1_c_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__1094),
            .in2(N__1181),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\generator_inst1.un3_counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.counter_2_LC_11_17_1 .C_ON=1'b1;
    defparam \generator_inst1.counter_2_LC_11_17_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_2_LC_11_17_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \generator_inst1.counter_2_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1239),
            .in3(N__619),
            .lcout(\generator_inst1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_1 ),
            .carryout(\generator_inst1.un3_counter_1_cry_2 ),
            .clk(N__1152),
            .ce(),
            .sr(N__1128));
    defparam \generator_inst1.counter_3_LC_11_17_2 .C_ON=1'b1;
    defparam \generator_inst1.counter_3_LC_11_17_2 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_3_LC_11_17_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \generator_inst1.counter_3_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1275),
            .in3(N__616),
            .lcout(\generator_inst1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_2 ),
            .carryout(\generator_inst1.un3_counter_1_cry_3 ),
            .clk(N__1152),
            .ce(),
            .sr(N__1128));
    defparam \generator_inst1.counter_4_LC_11_17_3 .C_ON=1'b1;
    defparam \generator_inst1.counter_4_LC_11_17_3 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_4_LC_11_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \generator_inst1.counter_4_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__1107),
            .in2(_gnd_net_),
            .in3(N__877),
            .lcout(\generator_inst1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_3 ),
            .carryout(\generator_inst1.un3_counter_1_cry_4 ),
            .clk(N__1152),
            .ce(),
            .sr(N__1128));
    defparam \generator_inst1.counter_5_LC_11_17_4 .C_ON=1'b1;
    defparam \generator_inst1.counter_5_LC_11_17_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_5_LC_11_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \generator_inst1.counter_5_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__873),
            .in2(_gnd_net_),
            .in3(N__862),
            .lcout(\generator_inst1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_4 ),
            .carryout(\generator_inst1.un3_counter_1_cry_5 ),
            .clk(N__1152),
            .ce(),
            .sr(N__1128));
    defparam \generator_inst1.counter_6_LC_11_17_5 .C_ON=1'b1;
    defparam \generator_inst1.counter_6_LC_11_17_5 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_6_LC_11_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \generator_inst1.counter_6_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__855),
            .in2(_gnd_net_),
            .in3(N__844),
            .lcout(\generator_inst1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_5 ),
            .carryout(\generator_inst1.un3_counter_1_cry_6 ),
            .clk(N__1152),
            .ce(),
            .sr(N__1128));
    defparam \generator_inst1.counter_7_LC_11_17_6 .C_ON=1'b1;
    defparam \generator_inst1.counter_7_LC_11_17_6 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_7_LC_11_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \generator_inst1.counter_7_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__840),
            .in2(_gnd_net_),
            .in3(N__829),
            .lcout(\generator_inst1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_6 ),
            .carryout(\generator_inst1.un3_counter_1_cry_7 ),
            .clk(N__1152),
            .ce(),
            .sr(N__1128));
    defparam \generator_inst1.counter_8_LC_11_17_7 .C_ON=1'b1;
    defparam \generator_inst1.counter_8_LC_11_17_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_8_LC_11_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \generator_inst1.counter_8_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__825),
            .in2(_gnd_net_),
            .in3(N__814),
            .lcout(\generator_inst1.counterZ0Z_8 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_7 ),
            .carryout(\generator_inst1.un3_counter_1_cry_8 ),
            .clk(N__1152),
            .ce(),
            .sr(N__1128));
    defparam \generator_inst1.counter_RNO_0_9_LC_11_18_0 .C_ON=1'b1;
    defparam \generator_inst1.counter_RNO_0_9_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.counter_RNO_0_9_LC_11_18_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \generator_inst1.counter_RNO_0_9_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__810),
            .in3(N__787),
            .lcout(\generator_inst1.counter_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\generator_inst1.un3_counter_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.counter_10_LC_11_18_1 .C_ON=1'b1;
    defparam \generator_inst1.counter_10_LC_11_18_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_10_LC_11_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \generator_inst1.counter_10_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__780),
            .in2(_gnd_net_),
            .in3(N__769),
            .lcout(\generator_inst1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_9 ),
            .carryout(\generator_inst1.un3_counter_1_cry_10 ),
            .clk(N__1155),
            .ce(),
            .sr(N__1130));
    defparam \generator_inst1.counter_11_LC_11_18_2 .C_ON=1'b1;
    defparam \generator_inst1.counter_11_LC_11_18_2 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_11_LC_11_18_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \generator_inst1.counter_11_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1293),
            .in3(N__766),
            .lcout(\generator_inst1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_10 ),
            .carryout(\generator_inst1.un3_counter_1_cry_11 ),
            .clk(N__1155),
            .ce(),
            .sr(N__1130));
    defparam \generator_inst1.counter_RNO_0_12_LC_11_18_3 .C_ON=1'b1;
    defparam \generator_inst1.counter_RNO_0_12_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.counter_RNO_0_12_LC_11_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \generator_inst1.counter_RNO_0_12_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__762),
            .in2(_gnd_net_),
            .in3(N__742),
            .lcout(\generator_inst1.counter_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_11 ),
            .carryout(\generator_inst1.un3_counter_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.counter_13_LC_11_18_4 .C_ON=1'b1;
    defparam \generator_inst1.counter_13_LC_11_18_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_13_LC_11_18_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \generator_inst1.counter_13_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__999),
            .in3(N__982),
            .lcout(\generator_inst1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_12 ),
            .carryout(\generator_inst1.un3_counter_1_cry_13 ),
            .clk(N__1155),
            .ce(),
            .sr(N__1130));
    defparam \generator_inst1.counter_14_LC_11_18_5 .C_ON=1'b1;
    defparam \generator_inst1.counter_14_LC_11_18_5 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_14_LC_11_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \generator_inst1.counter_14_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__1074),
            .in2(_gnd_net_),
            .in3(N__979),
            .lcout(\generator_inst1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_13 ),
            .carryout(\generator_inst1.un3_counter_1_cry_14 ),
            .clk(N__1155),
            .ce(),
            .sr(N__1130));
    defparam \generator_inst1.counter_15_LC_11_18_6 .C_ON=1'b1;
    defparam \generator_inst1.counter_15_LC_11_18_6 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_15_LC_11_18_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \generator_inst1.counter_15_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1063),
            .in3(N__976),
            .lcout(\generator_inst1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_14 ),
            .carryout(\generator_inst1.un3_counter_1_cry_15 ),
            .clk(N__1155),
            .ce(),
            .sr(N__1130));
    defparam \generator_inst1.counter_16_LC_11_18_7 .C_ON=1'b1;
    defparam \generator_inst1.counter_16_LC_11_18_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_16_LC_11_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \generator_inst1.counter_16_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(N__972),
            .in2(_gnd_net_),
            .in3(N__961),
            .lcout(\generator_inst1.counterZ0Z_16 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_15 ),
            .carryout(\generator_inst1.un3_counter_1_cry_16 ),
            .clk(N__1155),
            .ce(),
            .sr(N__1130));
    defparam \generator_inst1.counter_RNO_0_17_LC_11_19_0 .C_ON=1'b1;
    defparam \generator_inst1.counter_RNO_0_17_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.counter_RNO_0_17_LC_11_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \generator_inst1.counter_RNO_0_17_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__957),
            .in2(_gnd_net_),
            .in3(N__937),
            .lcout(\generator_inst1.counter_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\generator_inst1.un3_counter_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.counter_18_LC_11_19_1 .C_ON=1'b1;
    defparam \generator_inst1.counter_18_LC_11_19_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_18_LC_11_19_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \generator_inst1.counter_18_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1257),
            .in3(N__934),
            .lcout(\generator_inst1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_17 ),
            .carryout(\generator_inst1.un3_counter_1_cry_18 ),
            .clk(N__1156),
            .ce(),
            .sr(N__1132));
    defparam \generator_inst1.counter_RNO_0_19_LC_11_19_2 .C_ON=1'b1;
    defparam \generator_inst1.counter_RNO_0_19_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.counter_RNO_0_19_LC_11_19_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \generator_inst1.counter_RNO_0_19_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__931),
            .in3(N__907),
            .lcout(\generator_inst1.counter_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_18 ),
            .carryout(\generator_inst1.un3_counter_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.counter_RNO_0_20_LC_11_19_3 .C_ON=1'b1;
    defparam \generator_inst1.counter_RNO_0_20_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.counter_RNO_0_20_LC_11_19_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \generator_inst1.counter_RNO_0_20_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__903),
            .in3(N__880),
            .lcout(\generator_inst1.counter_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_19 ),
            .carryout(\generator_inst1.un3_counter_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.counter_RNO_0_21_LC_11_19_4 .C_ON=1'b1;
    defparam \generator_inst1.counter_RNO_0_21_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.counter_RNO_0_21_LC_11_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \generator_inst1.counter_RNO_0_21_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(N__1353),
            .in2(_gnd_net_),
            .in3(N__1336),
            .lcout(\generator_inst1.counter_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_20 ),
            .carryout(\generator_inst1.un3_counter_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.counter_RNO_0_22_LC_11_19_5 .C_ON=1'b1;
    defparam \generator_inst1.counter_RNO_0_22_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.counter_RNO_0_22_LC_11_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \generator_inst1.counter_RNO_0_22_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(N__1333),
            .in2(_gnd_net_),
            .in3(N__1315),
            .lcout(\generator_inst1.counter_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\generator_inst1.un3_counter_1_cry_21 ),
            .carryout(\generator_inst1.un3_counter_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.counter_23_LC_11_19_6 .C_ON=1'b0;
    defparam \generator_inst1.counter_23_LC_11_19_6 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_23_LC_11_19_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \generator_inst1.counter_23_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(N__1308),
            .in2(_gnd_net_),
            .in3(N__1312),
            .lcout(\generator_inst1.counterZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1156),
            .ce(),
            .sr(N__1132));
    defparam \generator_inst1.counter_RNISM7B1_2_LC_11_20_0 .C_ON=1'b0;
    defparam \generator_inst1.counter_RNISM7B1_2_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.counter_RNISM7B1_2_LC_11_20_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \generator_inst1.counter_RNISM7B1_2_LC_11_20_0  (
            .in0(N__1294),
            .in1(N__1276),
            .in2(N__1258),
            .in3(N__1240),
            .lcout(\generator_inst1.signal_out5_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.counter_1_LC_12_17_0 .C_ON=1'b0;
    defparam \generator_inst1.counter_1_LC_12_17_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.counter_1_LC_12_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \generator_inst1.counter_1_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__1182),
            .in2(_gnd_net_),
            .in3(N__1096),
            .lcout(\generator_inst1.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1153),
            .ce(),
            .sr(N__1131));
    defparam \generator_inst1.counter_RNISM7B1_1_LC_12_18_7 .C_ON=1'b0;
    defparam \generator_inst1.counter_RNISM7B1_1_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.counter_RNISM7B1_1_LC_12_18_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \generator_inst1.counter_RNISM7B1_1_LC_12_18_7  (
            .in0(N__1108),
            .in1(N__1095),
            .in2(N__1078),
            .in3(N__1062),
            .lcout(\generator_inst1.signal_out5_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RST_N_ibuf_RNIBJGC_LC_30_10_4.C_ON=1'b0;
    defparam RST_N_ibuf_RNIBJGC_LC_30_10_4.SEQ_MODE=4'b0000;
    defparam RST_N_ibuf_RNIBJGC_LC_30_10_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 RST_N_ibuf_RNIBJGC_LC_30_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1039),
            .lcout(RST_N_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
