-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 18 2025 08:30:48

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    generated_signal : out std_logic;
    RST_N : in std_logic;
    ENFIN : out std_logic;
    CLK : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__1656\ : std_logic;
signal \N__1655\ : std_logic;
signal \N__1654\ : std_logic;
signal \N__1645\ : std_logic;
signal \N__1644\ : std_logic;
signal \N__1643\ : std_logic;
signal \N__1636\ : std_logic;
signal \N__1635\ : std_logic;
signal \N__1634\ : std_logic;
signal \N__1627\ : std_logic;
signal \N__1626\ : std_logic;
signal \N__1625\ : std_logic;
signal \N__1608\ : std_logic;
signal \N__1605\ : std_logic;
signal \N__1602\ : std_logic;
signal \N__1601\ : std_logic;
signal \N__1600\ : std_logic;
signal \N__1595\ : std_logic;
signal \N__1592\ : std_logic;
signal \N__1587\ : std_logic;
signal \N__1584\ : std_logic;
signal \N__1583\ : std_logic;
signal \N__1580\ : std_logic;
signal \N__1577\ : std_logic;
signal \N__1572\ : std_logic;
signal \N__1569\ : std_logic;
signal \N__1568\ : std_logic;
signal \N__1567\ : std_logic;
signal \N__1564\ : std_logic;
signal \N__1559\ : std_logic;
signal \N__1556\ : std_logic;
signal \N__1551\ : std_logic;
signal \N__1548\ : std_logic;
signal \N__1547\ : std_logic;
signal \N__1544\ : std_logic;
signal \N__1541\ : std_logic;
signal \N__1538\ : std_logic;
signal \N__1533\ : std_logic;
signal \N__1530\ : std_logic;
signal \N__1527\ : std_logic;
signal \N__1526\ : std_logic;
signal \N__1523\ : std_logic;
signal \N__1520\ : std_logic;
signal \N__1515\ : std_logic;
signal \N__1512\ : std_logic;
signal \N__1509\ : std_logic;
signal \N__1508\ : std_logic;
signal \N__1505\ : std_logic;
signal \N__1502\ : std_logic;
signal \N__1497\ : std_logic;
signal \N__1496\ : std_logic;
signal \N__1495\ : std_logic;
signal \N__1494\ : std_logic;
signal \N__1493\ : std_logic;
signal \N__1492\ : std_logic;
signal \N__1491\ : std_logic;
signal \N__1490\ : std_logic;
signal \N__1489\ : std_logic;
signal \N__1488\ : std_logic;
signal \N__1487\ : std_logic;
signal \N__1464\ : std_logic;
signal \N__1461\ : std_logic;
signal \N__1458\ : std_logic;
signal \N__1457\ : std_logic;
signal \N__1456\ : std_logic;
signal \N__1455\ : std_logic;
signal \N__1454\ : std_logic;
signal \N__1453\ : std_logic;
signal \N__1452\ : std_logic;
signal \N__1437\ : std_logic;
signal \N__1434\ : std_logic;
signal \N__1431\ : std_logic;
signal \N__1430\ : std_logic;
signal \N__1429\ : std_logic;
signal \N__1428\ : std_logic;
signal \N__1425\ : std_logic;
signal \N__1422\ : std_logic;
signal \N__1421\ : std_logic;
signal \N__1418\ : std_logic;
signal \N__1415\ : std_logic;
signal \N__1412\ : std_logic;
signal \N__1409\ : std_logic;
signal \N__1406\ : std_logic;
signal \N__1395\ : std_logic;
signal \N__1394\ : std_logic;
signal \N__1393\ : std_logic;
signal \N__1392\ : std_logic;
signal \N__1391\ : std_logic;
signal \N__1390\ : std_logic;
signal \N__1389\ : std_logic;
signal \N__1388\ : std_logic;
signal \N__1379\ : std_logic;
signal \N__1370\ : std_logic;
signal \N__1365\ : std_logic;
signal \N__1364\ : std_logic;
signal \N__1361\ : std_logic;
signal \N__1358\ : std_logic;
signal \N__1355\ : std_logic;
signal \N__1350\ : std_logic;
signal \N__1347\ : std_logic;
signal \N__1344\ : std_logic;
signal \N__1343\ : std_logic;
signal \N__1338\ : std_logic;
signal \N__1335\ : std_logic;
signal \N__1334\ : std_logic;
signal \N__1333\ : std_logic;
signal \N__1332\ : std_logic;
signal \N__1331\ : std_logic;
signal \N__1330\ : std_logic;
signal \N__1329\ : std_logic;
signal \N__1328\ : std_logic;
signal \N__1327\ : std_logic;
signal \N__1326\ : std_logic;
signal \N__1323\ : std_logic;
signal \N__1320\ : std_logic;
signal \N__1317\ : std_logic;
signal \N__1314\ : std_logic;
signal \N__1305\ : std_logic;
signal \N__1300\ : std_logic;
signal \N__1287\ : std_logic;
signal \N__1286\ : std_logic;
signal \N__1283\ : std_logic;
signal \N__1280\ : std_logic;
signal \N__1277\ : std_logic;
signal \N__1274\ : std_logic;
signal \N__1269\ : std_logic;
signal \N__1268\ : std_logic;
signal \N__1267\ : std_logic;
signal \N__1264\ : std_logic;
signal \N__1263\ : std_logic;
signal \N__1260\ : std_logic;
signal \N__1257\ : std_logic;
signal \N__1254\ : std_logic;
signal \N__1251\ : std_logic;
signal \N__1248\ : std_logic;
signal \N__1245\ : std_logic;
signal \N__1240\ : std_logic;
signal \N__1235\ : std_logic;
signal \N__1232\ : std_logic;
signal \N__1229\ : std_logic;
signal \N__1224\ : std_logic;
signal \N__1223\ : std_logic;
signal \N__1222\ : std_logic;
signal \N__1221\ : std_logic;
signal \N__1220\ : std_logic;
signal \N__1219\ : std_logic;
signal \N__1218\ : std_logic;
signal \N__1217\ : std_logic;
signal \N__1216\ : std_logic;
signal \N__1215\ : std_logic;
signal \N__1214\ : std_logic;
signal \N__1213\ : std_logic;
signal \N__1212\ : std_logic;
signal \N__1211\ : std_logic;
signal \N__1210\ : std_logic;
signal \N__1207\ : std_logic;
signal \N__1206\ : std_logic;
signal \N__1205\ : std_logic;
signal \N__1202\ : std_logic;
signal \N__1187\ : std_logic;
signal \N__1174\ : std_logic;
signal \N__1171\ : std_logic;
signal \N__1166\ : std_logic;
signal \N__1155\ : std_logic;
signal \N__1154\ : std_logic;
signal \N__1151\ : std_logic;
signal \N__1148\ : std_logic;
signal \N__1143\ : std_logic;
signal \N__1140\ : std_logic;
signal \N__1137\ : std_logic;
signal \N__1134\ : std_logic;
signal \N__1133\ : std_logic;
signal \N__1132\ : std_logic;
signal \N__1127\ : std_logic;
signal \N__1124\ : std_logic;
signal \N__1119\ : std_logic;
signal \N__1116\ : std_logic;
signal \N__1113\ : std_logic;
signal \N__1112\ : std_logic;
signal \N__1111\ : std_logic;
signal \N__1108\ : std_logic;
signal \N__1105\ : std_logic;
signal \N__1102\ : std_logic;
signal \N__1095\ : std_logic;
signal \N__1092\ : std_logic;
signal \N__1089\ : std_logic;
signal \N__1086\ : std_logic;
signal \N__1083\ : std_logic;
signal \N__1080\ : std_logic;
signal \N__1077\ : std_logic;
signal \N__1074\ : std_logic;
signal \N__1071\ : std_logic;
signal \N__1068\ : std_logic;
signal \N__1065\ : std_logic;
signal \N__1062\ : std_logic;
signal \N__1059\ : std_logic;
signal \N__1056\ : std_logic;
signal \N__1053\ : std_logic;
signal \N__1050\ : std_logic;
signal \N__1047\ : std_logic;
signal \N__1046\ : std_logic;
signal \N__1045\ : std_logic;
signal \N__1044\ : std_logic;
signal \N__1041\ : std_logic;
signal \N__1040\ : std_logic;
signal \N__1039\ : std_logic;
signal \N__1036\ : std_logic;
signal \N__1027\ : std_logic;
signal \N__1024\ : std_logic;
signal \N__1017\ : std_logic;
signal \N__1014\ : std_logic;
signal \N__1011\ : std_logic;
signal \N__1010\ : std_logic;
signal \N__1009\ : std_logic;
signal \N__1008\ : std_logic;
signal \N__1005\ : std_logic;
signal \N__1002\ : std_logic;
signal \N__1001\ : std_logic;
signal \N__996\ : std_logic;
signal \N__989\ : std_logic;
signal \N__984\ : std_logic;
signal \N__983\ : std_logic;
signal \N__982\ : std_logic;
signal \N__981\ : std_logic;
signal \N__980\ : std_logic;
signal \N__977\ : std_logic;
signal \N__976\ : std_logic;
signal \N__973\ : std_logic;
signal \N__970\ : std_logic;
signal \N__961\ : std_logic;
signal \N__954\ : std_logic;
signal \N__953\ : std_logic;
signal \N__952\ : std_logic;
signal \N__951\ : std_logic;
signal \N__950\ : std_logic;
signal \N__947\ : std_logic;
signal \N__944\ : std_logic;
signal \N__937\ : std_logic;
signal \N__934\ : std_logic;
signal \N__927\ : std_logic;
signal \N__924\ : std_logic;
signal \N__923\ : std_logic;
signal \N__922\ : std_logic;
signal \N__921\ : std_logic;
signal \N__918\ : std_logic;
signal \N__911\ : std_logic;
signal \N__906\ : std_logic;
signal \N__903\ : std_logic;
signal \N__900\ : std_logic;
signal \N__897\ : std_logic;
signal \N__894\ : std_logic;
signal \N__891\ : std_logic;
signal \N__888\ : std_logic;
signal \N__885\ : std_logic;
signal \N__882\ : std_logic;
signal \N__879\ : std_logic;
signal \N__876\ : std_logic;
signal \N__873\ : std_logic;
signal \N__870\ : std_logic;
signal \N__867\ : std_logic;
signal \N__864\ : std_logic;
signal \N__861\ : std_logic;
signal \N__858\ : std_logic;
signal \N__857\ : std_logic;
signal \N__856\ : std_logic;
signal \N__855\ : std_logic;
signal \N__854\ : std_logic;
signal \N__851\ : std_logic;
signal \N__842\ : std_logic;
signal \N__837\ : std_logic;
signal \N__836\ : std_logic;
signal \N__835\ : std_logic;
signal \N__834\ : std_logic;
signal \N__831\ : std_logic;
signal \N__824\ : std_logic;
signal \N__819\ : std_logic;
signal \N__816\ : std_logic;
signal \N__815\ : std_logic;
signal \N__814\ : std_logic;
signal \N__813\ : std_logic;
signal \N__810\ : std_logic;
signal \N__803\ : std_logic;
signal \N__798\ : std_logic;
signal \N__795\ : std_logic;
signal \N__792\ : std_logic;
signal \N__789\ : std_logic;
signal \N__786\ : std_logic;
signal \N__783\ : std_logic;
signal \N__780\ : std_logic;
signal \N__779\ : std_logic;
signal \N__776\ : std_logic;
signal \N__775\ : std_logic;
signal \N__768\ : std_logic;
signal \N__765\ : std_logic;
signal \N__762\ : std_logic;
signal \N__759\ : std_logic;
signal \N__758\ : std_logic;
signal \N__755\ : std_logic;
signal \N__752\ : std_logic;
signal \N__747\ : std_logic;
signal \N__744\ : std_logic;
signal \N__741\ : std_logic;
signal \N__738\ : std_logic;
signal \N__735\ : std_logic;
signal \N__732\ : std_logic;
signal \N__729\ : std_logic;
signal \N__726\ : std_logic;
signal \N__723\ : std_logic;
signal \N__720\ : std_logic;
signal \N__717\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal signal_out_fsm : std_logic;
signal \SELSTAT\ : std_logic;
signal \SELDYN\ : std_logic;
signal generated_signal_c : std_logic;
signal \RST_N_c_i\ : std_logic;
signal \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.N_125_1_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.counterZ0Z_0\ : std_logic;
signal \fsm_shiftRegs_inst1.counterZ0Z_1\ : std_logic;
signal \fsm_shiftRegs_inst1.counterZ0Z_2\ : std_logic;
signal \fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.N_125_1\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2\ : std_logic;
signal \fsm_shiftRegs_inst1.counterDYNZ0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.counterDYNZ0Z_2\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_15\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_14\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_13\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_12\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_11\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_10\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_5\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_6\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_4\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_7\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_8\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_9\ : std_logic;
signal \ENFIN_c\ : std_logic;
signal \fsm_shiftRegs_inst1.current_stateZ0Z_1\ : std_logic;
signal \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.counterZ0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.counterDYNZ0Z_0\ : std_logic;
signal \fsm_shiftRegs_inst1.counterDYNZ0Z_1\ : std_logic;
signal \fsm_shiftRegs_inst1.current_stateZ0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0\ : std_logic;
signal \fsm_shiftRegs_inst1.current_stateZ0Z_2\ : std_logic;
signal \fsm_shiftRegs_inst1.un1_current_state4_0\ : std_logic;
signal \RST_N_c\ : std_logic;
signal \fsm_shiftRegs_inst1.current_stateZ0Z_0\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_2\ : std_logic;
signal \fsm_shiftRegs_inst1.N_122_i\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_0\ : std_logic;
signal \bfn_4_11_0_\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_1\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_0\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_2\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_1\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_2\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_4\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_3\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_5\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_4\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_6\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_5\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_6\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_7\ : std_logic;
signal \CLK_c_g\ : std_logic;
signal \RST_N_c_i_g\ : std_logic;
signal \fsm_shiftRegs_inst1.current_stateZ0Z_4\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_i_4\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \RST_N_wire\ : std_logic;
signal \ENFIN_wire\ : std_logic;
signal generated_signal_wire : std_logic;

begin
    \CLK_wire\ <= CLK;
    \RST_N_wire\ <= RST_N;
    ENFIN <= \ENFIN_wire\;
    generated_signal <= generated_signal_wire;

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__1654\,
            GLOBALBUFFEROUTPUT => \CLK_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1656\,
            DIN => \N__1655\,
            DOUT => \N__1654\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1656\,
            PADOUT => \N__1655\,
            PADIN => \N__1654\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RST_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1645\,
            DIN => \N__1644\,
            DOUT => \N__1643\,
            PACKAGEPIN => \RST_N_wire\
        );

    \RST_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1645\,
            PADOUT => \N__1644\,
            PADIN => \N__1643\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RST_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ENFIN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1636\,
            DIN => \N__1635\,
            DOUT => \N__1634\,
            PACKAGEPIN => \ENFIN_wire\
        );

    \ENFIN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1636\,
            PADOUT => \N__1635\,
            PADIN => \N__1634\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1059\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \generated_signal_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1627\,
            DIN => \N__1626\,
            DOUT => \N__1625\,
            PACKAGEPIN => generated_signal_wire
        );

    \generated_signal_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1627\,
            PADOUT => \N__1626\,
            PADIN => \N__1625\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__735\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__360\ : InMux
    port map (
            O => \N__1608\,
            I => \fsm_shiftRegs_inst1.counter2_cry_0\
        );

    \I__359\ : CascadeMux
    port map (
            O => \N__1605\,
            I => \N__1602\
        );

    \I__358\ : InMux
    port map (
            O => \N__1602\,
            I => \N__1595\
        );

    \I__357\ : InMux
    port map (
            O => \N__1601\,
            I => \N__1595\
        );

    \I__356\ : InMux
    port map (
            O => \N__1600\,
            I => \N__1592\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__1595\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_2\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__1592\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_2\
        );

    \I__353\ : InMux
    port map (
            O => \N__1587\,
            I => \fsm_shiftRegs_inst1.counter2_cry_1\
        );

    \I__352\ : InMux
    port map (
            O => \N__1584\,
            I => \N__1580\
        );

    \I__351\ : InMux
    port map (
            O => \N__1583\,
            I => \N__1577\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__1580\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_3\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__1577\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_3\
        );

    \I__348\ : InMux
    port map (
            O => \N__1572\,
            I => \fsm_shiftRegs_inst1.counter2_cry_2\
        );

    \I__347\ : CascadeMux
    port map (
            O => \N__1569\,
            I => \N__1564\
        );

    \I__346\ : InMux
    port map (
            O => \N__1568\,
            I => \N__1559\
        );

    \I__345\ : InMux
    port map (
            O => \N__1567\,
            I => \N__1559\
        );

    \I__344\ : InMux
    port map (
            O => \N__1564\,
            I => \N__1556\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__1559\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_4\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__1556\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_4\
        );

    \I__341\ : InMux
    port map (
            O => \N__1551\,
            I => \fsm_shiftRegs_inst1.counter2_cry_3\
        );

    \I__340\ : CascadeMux
    port map (
            O => \N__1548\,
            I => \N__1544\
        );

    \I__339\ : InMux
    port map (
            O => \N__1547\,
            I => \N__1541\
        );

    \I__338\ : InMux
    port map (
            O => \N__1544\,
            I => \N__1538\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__1541\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_5\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__1538\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_5\
        );

    \I__335\ : InMux
    port map (
            O => \N__1533\,
            I => \fsm_shiftRegs_inst1.counter2_cry_4\
        );

    \I__334\ : CascadeMux
    port map (
            O => \N__1530\,
            I => \N__1527\
        );

    \I__333\ : InMux
    port map (
            O => \N__1527\,
            I => \N__1523\
        );

    \I__332\ : InMux
    port map (
            O => \N__1526\,
            I => \N__1520\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__1523\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_6\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__1520\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_6\
        );

    \I__329\ : InMux
    port map (
            O => \N__1515\,
            I => \fsm_shiftRegs_inst1.counter2_cry_5\
        );

    \I__328\ : InMux
    port map (
            O => \N__1512\,
            I => \fsm_shiftRegs_inst1.counter2_cry_6\
        );

    \I__327\ : InMux
    port map (
            O => \N__1509\,
            I => \N__1505\
        );

    \I__326\ : InMux
    port map (
            O => \N__1508\,
            I => \N__1502\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__1505\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_7\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__1502\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_7\
        );

    \I__323\ : ClkMux
    port map (
            O => \N__1497\,
            I => \N__1464\
        );

    \I__322\ : ClkMux
    port map (
            O => \N__1496\,
            I => \N__1464\
        );

    \I__321\ : ClkMux
    port map (
            O => \N__1495\,
            I => \N__1464\
        );

    \I__320\ : ClkMux
    port map (
            O => \N__1494\,
            I => \N__1464\
        );

    \I__319\ : ClkMux
    port map (
            O => \N__1493\,
            I => \N__1464\
        );

    \I__318\ : ClkMux
    port map (
            O => \N__1492\,
            I => \N__1464\
        );

    \I__317\ : ClkMux
    port map (
            O => \N__1491\,
            I => \N__1464\
        );

    \I__316\ : ClkMux
    port map (
            O => \N__1490\,
            I => \N__1464\
        );

    \I__315\ : ClkMux
    port map (
            O => \N__1489\,
            I => \N__1464\
        );

    \I__314\ : ClkMux
    port map (
            O => \N__1488\,
            I => \N__1464\
        );

    \I__313\ : ClkMux
    port map (
            O => \N__1487\,
            I => \N__1464\
        );

    \I__312\ : GlobalMux
    port map (
            O => \N__1464\,
            I => \N__1461\
        );

    \I__311\ : gio2CtrlBuf
    port map (
            O => \N__1461\,
            I => \CLK_c_g\
        );

    \I__310\ : SRMux
    port map (
            O => \N__1458\,
            I => \N__1437\
        );

    \I__309\ : SRMux
    port map (
            O => \N__1457\,
            I => \N__1437\
        );

    \I__308\ : SRMux
    port map (
            O => \N__1456\,
            I => \N__1437\
        );

    \I__307\ : SRMux
    port map (
            O => \N__1455\,
            I => \N__1437\
        );

    \I__306\ : SRMux
    port map (
            O => \N__1454\,
            I => \N__1437\
        );

    \I__305\ : SRMux
    port map (
            O => \N__1453\,
            I => \N__1437\
        );

    \I__304\ : SRMux
    port map (
            O => \N__1452\,
            I => \N__1437\
        );

    \I__303\ : GlobalMux
    port map (
            O => \N__1437\,
            I => \N__1434\
        );

    \I__302\ : gio2CtrlBuf
    port map (
            O => \N__1434\,
            I => \RST_N_c_i_g\
        );

    \I__301\ : InMux
    port map (
            O => \N__1431\,
            I => \N__1425\
        );

    \I__300\ : InMux
    port map (
            O => \N__1430\,
            I => \N__1422\
        );

    \I__299\ : InMux
    port map (
            O => \N__1429\,
            I => \N__1418\
        );

    \I__298\ : InMux
    port map (
            O => \N__1428\,
            I => \N__1415\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__1425\,
            I => \N__1412\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__1422\,
            I => \N__1409\
        );

    \I__295\ : InMux
    port map (
            O => \N__1421\,
            I => \N__1406\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__1418\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_4\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__1415\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_4\
        );

    \I__292\ : Odrv4
    port map (
            O => \N__1412\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_4\
        );

    \I__291\ : Odrv4
    port map (
            O => \N__1409\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_4\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__1406\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_4\
        );

    \I__289\ : InMux
    port map (
            O => \N__1395\,
            I => \N__1379\
        );

    \I__288\ : InMux
    port map (
            O => \N__1394\,
            I => \N__1379\
        );

    \I__287\ : InMux
    port map (
            O => \N__1393\,
            I => \N__1379\
        );

    \I__286\ : InMux
    port map (
            O => \N__1392\,
            I => \N__1379\
        );

    \I__285\ : InMux
    port map (
            O => \N__1391\,
            I => \N__1370\
        );

    \I__284\ : InMux
    port map (
            O => \N__1390\,
            I => \N__1370\
        );

    \I__283\ : InMux
    port map (
            O => \N__1389\,
            I => \N__1370\
        );

    \I__282\ : InMux
    port map (
            O => \N__1388\,
            I => \N__1370\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__1379\,
            I => \fsm_shiftRegs_inst1.current_state_i_4\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__1370\,
            I => \fsm_shiftRegs_inst1.current_state_i_4\
        );

    \I__279\ : InMux
    port map (
            O => \N__1365\,
            I => \N__1361\
        );

    \I__278\ : InMux
    port map (
            O => \N__1364\,
            I => \N__1358\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__1361\,
            I => \N__1355\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__1358\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_3\
        );

    \I__275\ : Odrv12
    port map (
            O => \N__1355\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_3\
        );

    \I__274\ : CascadeMux
    port map (
            O => \N__1350\,
            I => \fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_\
        );

    \I__273\ : CascadeMux
    port map (
            O => \N__1347\,
            I => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_\
        );

    \I__272\ : InMux
    port map (
            O => \N__1344\,
            I => \N__1338\
        );

    \I__271\ : InMux
    port map (
            O => \N__1343\,
            I => \N__1338\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__1338\,
            I => \fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0\
        );

    \I__269\ : InMux
    port map (
            O => \N__1335\,
            I => \N__1323\
        );

    \I__268\ : InMux
    port map (
            O => \N__1334\,
            I => \N__1320\
        );

    \I__267\ : InMux
    port map (
            O => \N__1333\,
            I => \N__1317\
        );

    \I__266\ : InMux
    port map (
            O => \N__1332\,
            I => \N__1314\
        );

    \I__265\ : InMux
    port map (
            O => \N__1331\,
            I => \N__1305\
        );

    \I__264\ : InMux
    port map (
            O => \N__1330\,
            I => \N__1305\
        );

    \I__263\ : InMux
    port map (
            O => \N__1329\,
            I => \N__1305\
        );

    \I__262\ : InMux
    port map (
            O => \N__1328\,
            I => \N__1305\
        );

    \I__261\ : InMux
    port map (
            O => \N__1327\,
            I => \N__1300\
        );

    \I__260\ : InMux
    port map (
            O => \N__1326\,
            I => \N__1300\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__1323\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_2\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__1320\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_2\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__1317\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_2\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__1314\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_2\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__1305\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_2\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__1300\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_2\
        );

    \I__253\ : CEMux
    port map (
            O => \N__1287\,
            I => \N__1283\
        );

    \I__252\ : CEMux
    port map (
            O => \N__1286\,
            I => \N__1280\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__1283\,
            I => \N__1277\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__1280\,
            I => \N__1274\
        );

    \I__249\ : Odrv4
    port map (
            O => \N__1277\,
            I => \fsm_shiftRegs_inst1.un1_current_state4_0\
        );

    \I__248\ : Odrv4
    port map (
            O => \N__1274\,
            I => \fsm_shiftRegs_inst1.un1_current_state4_0\
        );

    \I__247\ : InMux
    port map (
            O => \N__1269\,
            I => \N__1264\
        );

    \I__246\ : InMux
    port map (
            O => \N__1268\,
            I => \N__1260\
        );

    \I__245\ : CascadeMux
    port map (
            O => \N__1267\,
            I => \N__1257\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__1264\,
            I => \N__1254\
        );

    \I__243\ : InMux
    port map (
            O => \N__1263\,
            I => \N__1251\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__1260\,
            I => \N__1248\
        );

    \I__241\ : InMux
    port map (
            O => \N__1257\,
            I => \N__1245\
        );

    \I__240\ : Span4Mux_v
    port map (
            O => \N__1254\,
            I => \N__1240\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__1251\,
            I => \N__1240\
        );

    \I__238\ : Span4Mux_v
    port map (
            O => \N__1248\,
            I => \N__1235\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__1245\,
            I => \N__1235\
        );

    \I__236\ : Span4Mux_v
    port map (
            O => \N__1240\,
            I => \N__1232\
        );

    \I__235\ : Span4Mux_v
    port map (
            O => \N__1235\,
            I => \N__1229\
        );

    \I__234\ : Odrv4
    port map (
            O => \N__1232\,
            I => \RST_N_c\
        );

    \I__233\ : Odrv4
    port map (
            O => \N__1229\,
            I => \RST_N_c\
        );

    \I__232\ : InMux
    port map (
            O => \N__1224\,
            I => \N__1207\
        );

    \I__231\ : InMux
    port map (
            O => \N__1223\,
            I => \N__1202\
        );

    \I__230\ : InMux
    port map (
            O => \N__1222\,
            I => \N__1187\
        );

    \I__229\ : InMux
    port map (
            O => \N__1221\,
            I => \N__1187\
        );

    \I__228\ : InMux
    port map (
            O => \N__1220\,
            I => \N__1187\
        );

    \I__227\ : InMux
    port map (
            O => \N__1219\,
            I => \N__1187\
        );

    \I__226\ : InMux
    port map (
            O => \N__1218\,
            I => \N__1187\
        );

    \I__225\ : InMux
    port map (
            O => \N__1217\,
            I => \N__1187\
        );

    \I__224\ : InMux
    port map (
            O => \N__1216\,
            I => \N__1187\
        );

    \I__223\ : InMux
    port map (
            O => \N__1215\,
            I => \N__1174\
        );

    \I__222\ : InMux
    port map (
            O => \N__1214\,
            I => \N__1174\
        );

    \I__221\ : InMux
    port map (
            O => \N__1213\,
            I => \N__1174\
        );

    \I__220\ : InMux
    port map (
            O => \N__1212\,
            I => \N__1174\
        );

    \I__219\ : InMux
    port map (
            O => \N__1211\,
            I => \N__1174\
        );

    \I__218\ : InMux
    port map (
            O => \N__1210\,
            I => \N__1174\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__1207\,
            I => \N__1171\
        );

    \I__216\ : InMux
    port map (
            O => \N__1206\,
            I => \N__1166\
        );

    \I__215\ : InMux
    port map (
            O => \N__1205\,
            I => \N__1166\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__1202\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_0\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__1187\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_0\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__1174\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_0\
        );

    \I__211\ : Odrv4
    port map (
            O => \N__1171\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_0\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__1166\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_0\
        );

    \I__209\ : InMux
    port map (
            O => \N__1155\,
            I => \N__1151\
        );

    \I__208\ : InMux
    port map (
            O => \N__1154\,
            I => \N__1148\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__1151\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_2\
        );

    \I__206\ : LocalMux
    port map (
            O => \N__1148\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_2\
        );

    \I__205\ : CEMux
    port map (
            O => \N__1143\,
            I => \N__1140\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__1140\,
            I => \N__1137\
        );

    \I__203\ : Odrv12
    port map (
            O => \N__1137\,
            I => \fsm_shiftRegs_inst1.N_122_i\
        );

    \I__202\ : InMux
    port map (
            O => \N__1134\,
            I => \N__1127\
        );

    \I__201\ : InMux
    port map (
            O => \N__1133\,
            I => \N__1127\
        );

    \I__200\ : InMux
    port map (
            O => \N__1132\,
            I => \N__1124\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__1127\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_0\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__1124\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_0\
        );

    \I__197\ : InMux
    port map (
            O => \N__1119\,
            I => \bfn_4_11_0_\
        );

    \I__196\ : InMux
    port map (
            O => \N__1116\,
            I => \N__1113\
        );

    \I__195\ : LocalMux
    port map (
            O => \N__1113\,
            I => \N__1108\
        );

    \I__194\ : InMux
    port map (
            O => \N__1112\,
            I => \N__1105\
        );

    \I__193\ : InMux
    port map (
            O => \N__1111\,
            I => \N__1102\
        );

    \I__192\ : Odrv4
    port map (
            O => \N__1108\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_1\
        );

    \I__191\ : LocalMux
    port map (
            O => \N__1105\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_1\
        );

    \I__190\ : LocalMux
    port map (
            O => \N__1102\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_1\
        );

    \I__189\ : InMux
    port map (
            O => \N__1095\,
            I => \N__1092\
        );

    \I__188\ : LocalMux
    port map (
            O => \N__1092\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_6\
        );

    \I__187\ : InMux
    port map (
            O => \N__1089\,
            I => \N__1086\
        );

    \I__186\ : LocalMux
    port map (
            O => \N__1086\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_3\
        );

    \I__185\ : InMux
    port map (
            O => \N__1083\,
            I => \N__1080\
        );

    \I__184\ : LocalMux
    port map (
            O => \N__1080\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_4\
        );

    \I__183\ : InMux
    port map (
            O => \N__1077\,
            I => \N__1074\
        );

    \I__182\ : LocalMux
    port map (
            O => \N__1074\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_7\
        );

    \I__181\ : InMux
    port map (
            O => \N__1071\,
            I => \N__1068\
        );

    \I__180\ : LocalMux
    port map (
            O => \N__1068\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_8\
        );

    \I__179\ : InMux
    port map (
            O => \N__1065\,
            I => \N__1062\
        );

    \I__178\ : LocalMux
    port map (
            O => \N__1062\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_9\
        );

    \I__177\ : IoInMux
    port map (
            O => \N__1059\,
            I => \N__1056\
        );

    \I__176\ : LocalMux
    port map (
            O => \N__1056\,
            I => \N__1053\
        );

    \I__175\ : Span4Mux_s1_h
    port map (
            O => \N__1053\,
            I => \N__1050\
        );

    \I__174\ : Odrv4
    port map (
            O => \N__1050\,
            I => \ENFIN_c\
        );

    \I__173\ : CascadeMux
    port map (
            O => \N__1047\,
            I => \N__1041\
        );

    \I__172\ : InMux
    port map (
            O => \N__1046\,
            I => \N__1036\
        );

    \I__171\ : InMux
    port map (
            O => \N__1045\,
            I => \N__1027\
        );

    \I__170\ : InMux
    port map (
            O => \N__1044\,
            I => \N__1027\
        );

    \I__169\ : InMux
    port map (
            O => \N__1041\,
            I => \N__1027\
        );

    \I__168\ : InMux
    port map (
            O => \N__1040\,
            I => \N__1027\
        );

    \I__167\ : InMux
    port map (
            O => \N__1039\,
            I => \N__1024\
        );

    \I__166\ : LocalMux
    port map (
            O => \N__1036\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_1\
        );

    \I__165\ : LocalMux
    port map (
            O => \N__1027\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_1\
        );

    \I__164\ : LocalMux
    port map (
            O => \N__1024\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_1\
        );

    \I__163\ : InMux
    port map (
            O => \N__1017\,
            I => \N__1014\
        );

    \I__162\ : LocalMux
    port map (
            O => \N__1014\,
            I => \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3\
        );

    \I__161\ : CascadeMux
    port map (
            O => \N__1011\,
            I => \N__1005\
        );

    \I__160\ : CascadeMux
    port map (
            O => \N__1010\,
            I => \N__1002\
        );

    \I__159\ : InMux
    port map (
            O => \N__1009\,
            I => \N__996\
        );

    \I__158\ : InMux
    port map (
            O => \N__1008\,
            I => \N__996\
        );

    \I__157\ : InMux
    port map (
            O => \N__1005\,
            I => \N__989\
        );

    \I__156\ : InMux
    port map (
            O => \N__1002\,
            I => \N__989\
        );

    \I__155\ : InMux
    port map (
            O => \N__1001\,
            I => \N__989\
        );

    \I__154\ : LocalMux
    port map (
            O => \N__996\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_3\
        );

    \I__153\ : LocalMux
    port map (
            O => \N__989\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_3\
        );

    \I__152\ : CascadeMux
    port map (
            O => \N__984\,
            I => \N__977\
        );

    \I__151\ : InMux
    port map (
            O => \N__983\,
            I => \N__973\
        );

    \I__150\ : InMux
    port map (
            O => \N__982\,
            I => \N__970\
        );

    \I__149\ : InMux
    port map (
            O => \N__981\,
            I => \N__961\
        );

    \I__148\ : InMux
    port map (
            O => \N__980\,
            I => \N__961\
        );

    \I__147\ : InMux
    port map (
            O => \N__977\,
            I => \N__961\
        );

    \I__146\ : InMux
    port map (
            O => \N__976\,
            I => \N__961\
        );

    \I__145\ : LocalMux
    port map (
            O => \N__973\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_0\
        );

    \I__144\ : LocalMux
    port map (
            O => \N__970\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_0\
        );

    \I__143\ : LocalMux
    port map (
            O => \N__961\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_0\
        );

    \I__142\ : CascadeMux
    port map (
            O => \N__954\,
            I => \N__947\
        );

    \I__141\ : InMux
    port map (
            O => \N__953\,
            I => \N__944\
        );

    \I__140\ : InMux
    port map (
            O => \N__952\,
            I => \N__937\
        );

    \I__139\ : InMux
    port map (
            O => \N__951\,
            I => \N__937\
        );

    \I__138\ : InMux
    port map (
            O => \N__950\,
            I => \N__937\
        );

    \I__137\ : InMux
    port map (
            O => \N__947\,
            I => \N__934\
        );

    \I__136\ : LocalMux
    port map (
            O => \N__944\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_1\
        );

    \I__135\ : LocalMux
    port map (
            O => \N__937\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_1\
        );

    \I__134\ : LocalMux
    port map (
            O => \N__934\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_1\
        );

    \I__133\ : CascadeMux
    port map (
            O => \N__927\,
            I => \N__924\
        );

    \I__132\ : InMux
    port map (
            O => \N__924\,
            I => \N__918\
        );

    \I__131\ : InMux
    port map (
            O => \N__923\,
            I => \N__911\
        );

    \I__130\ : InMux
    port map (
            O => \N__922\,
            I => \N__911\
        );

    \I__129\ : InMux
    port map (
            O => \N__921\,
            I => \N__911\
        );

    \I__128\ : LocalMux
    port map (
            O => \N__918\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_2\
        );

    \I__127\ : LocalMux
    port map (
            O => \N__911\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_2\
        );

    \I__126\ : InMux
    port map (
            O => \N__906\,
            I => \N__903\
        );

    \I__125\ : LocalMux
    port map (
            O => \N__903\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_15\
        );

    \I__124\ : InMux
    port map (
            O => \N__900\,
            I => \N__897\
        );

    \I__123\ : LocalMux
    port map (
            O => \N__897\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_14\
        );

    \I__122\ : InMux
    port map (
            O => \N__894\,
            I => \N__891\
        );

    \I__121\ : LocalMux
    port map (
            O => \N__891\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_13\
        );

    \I__120\ : InMux
    port map (
            O => \N__888\,
            I => \N__885\
        );

    \I__119\ : LocalMux
    port map (
            O => \N__885\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_12\
        );

    \I__118\ : InMux
    port map (
            O => \N__882\,
            I => \N__879\
        );

    \I__117\ : LocalMux
    port map (
            O => \N__879\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_11\
        );

    \I__116\ : InMux
    port map (
            O => \N__876\,
            I => \N__873\
        );

    \I__115\ : LocalMux
    port map (
            O => \N__873\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_10\
        );

    \I__114\ : InMux
    port map (
            O => \N__870\,
            I => \N__867\
        );

    \I__113\ : LocalMux
    port map (
            O => \N__867\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_5\
        );

    \I__112\ : CascadeMux
    port map (
            O => \N__864\,
            I => \fsm_shiftRegs_inst1.N_125_1_cascade_\
        );

    \I__111\ : CascadeMux
    port map (
            O => \N__861\,
            I => \N__858\
        );

    \I__110\ : InMux
    port map (
            O => \N__858\,
            I => \N__851\
        );

    \I__109\ : InMux
    port map (
            O => \N__857\,
            I => \N__842\
        );

    \I__108\ : InMux
    port map (
            O => \N__856\,
            I => \N__842\
        );

    \I__107\ : InMux
    port map (
            O => \N__855\,
            I => \N__842\
        );

    \I__106\ : InMux
    port map (
            O => \N__854\,
            I => \N__842\
        );

    \I__105\ : LocalMux
    port map (
            O => \N__851\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_0\
        );

    \I__104\ : LocalMux
    port map (
            O => \N__842\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_0\
        );

    \I__103\ : InMux
    port map (
            O => \N__837\,
            I => \N__831\
        );

    \I__102\ : InMux
    port map (
            O => \N__836\,
            I => \N__824\
        );

    \I__101\ : InMux
    port map (
            O => \N__835\,
            I => \N__824\
        );

    \I__100\ : InMux
    port map (
            O => \N__834\,
            I => \N__824\
        );

    \I__99\ : LocalMux
    port map (
            O => \N__831\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_1\
        );

    \I__98\ : LocalMux
    port map (
            O => \N__824\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_1\
        );

    \I__97\ : CascadeMux
    port map (
            O => \N__819\,
            I => \N__816\
        );

    \I__96\ : InMux
    port map (
            O => \N__816\,
            I => \N__810\
        );

    \I__95\ : InMux
    port map (
            O => \N__815\,
            I => \N__803\
        );

    \I__94\ : InMux
    port map (
            O => \N__814\,
            I => \N__803\
        );

    \I__93\ : InMux
    port map (
            O => \N__813\,
            I => \N__803\
        );

    \I__92\ : LocalMux
    port map (
            O => \N__810\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_2\
        );

    \I__91\ : LocalMux
    port map (
            O => \N__803\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_2\
        );

    \I__90\ : CascadeMux
    port map (
            O => \N__798\,
            I => \fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_\
        );

    \I__89\ : InMux
    port map (
            O => \N__795\,
            I => \N__792\
        );

    \I__88\ : LocalMux
    port map (
            O => \N__792\,
            I => \fsm_shiftRegs_inst1.N_125_1\
        );

    \I__87\ : CascadeMux
    port map (
            O => \N__789\,
            I => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_\
        );

    \I__86\ : InMux
    port map (
            O => \N__786\,
            I => \N__783\
        );

    \I__85\ : LocalMux
    port map (
            O => \N__783\,
            I => \fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2\
        );

    \I__84\ : CascadeMux
    port map (
            O => \N__780\,
            I => \N__776\
        );

    \I__83\ : InMux
    port map (
            O => \N__779\,
            I => \N__768\
        );

    \I__82\ : InMux
    port map (
            O => \N__776\,
            I => \N__768\
        );

    \I__81\ : InMux
    port map (
            O => \N__775\,
            I => \N__768\
        );

    \I__80\ : LocalMux
    port map (
            O => \N__768\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_3\
        );

    \I__79\ : InMux
    port map (
            O => \N__765\,
            I => \N__762\
        );

    \I__78\ : LocalMux
    port map (
            O => \N__762\,
            I => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3\
        );

    \I__77\ : InMux
    port map (
            O => \N__759\,
            I => \N__755\
        );

    \I__76\ : InMux
    port map (
            O => \N__758\,
            I => \N__752\
        );

    \I__75\ : LocalMux
    port map (
            O => \N__755\,
            I => signal_out_fsm
        );

    \I__74\ : LocalMux
    port map (
            O => \N__752\,
            I => signal_out_fsm
        );

    \I__73\ : InMux
    port map (
            O => \N__747\,
            I => \N__744\
        );

    \I__72\ : LocalMux
    port map (
            O => \N__744\,
            I => \SELSTAT\
        );

    \I__71\ : InMux
    port map (
            O => \N__741\,
            I => \N__738\
        );

    \I__70\ : LocalMux
    port map (
            O => \N__738\,
            I => \SELDYN\
        );

    \I__69\ : IoInMux
    port map (
            O => \N__735\,
            I => \N__732\
        );

    \I__68\ : LocalMux
    port map (
            O => \N__732\,
            I => \N__729\
        );

    \I__67\ : Span12Mux_s0_h
    port map (
            O => \N__729\,
            I => \N__726\
        );

    \I__66\ : Odrv12
    port map (
            O => \N__726\,
            I => generated_signal_c
        );

    \I__65\ : IoInMux
    port map (
            O => \N__723\,
            I => \N__720\
        );

    \I__64\ : LocalMux
    port map (
            O => \N__720\,
            I => \RST_N_c_i\
        );

    \I__63\ : CascadeMux
    port map (
            O => \N__717\,
            I => \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_\
        );

    \IN_MUX_bfv_4_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_11_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \RST_N_ibuf_RNIBJGC_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__723\,
            GLOBALBUFFEROUTPUT => \RST_N_c_i_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.signal_out_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__759\,
            in1 => \N__906\,
            in2 => \N__1267\,
            in3 => \N__1335\,
            lcout => signal_out_fsm,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_RNO_1_2_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__819\,
            in3 => \N__1039\,
            lcout => \fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.sel_stat_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1364\,
            lcout => \SELSTAT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1488\,
            ce => 'H',
            sr => \N__1453\
        );

    \fsm_shiftRegs_inst1.sel_dyn_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1333\,
            in2 => \_gnd_net_\,
            in3 => \N__1431\,
            lcout => \SELDYN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1488\,
            ce => 'H',
            sr => \N__1453\
        );

    \generator_inst1.signal_aux_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__758\,
            in1 => \N__747\,
            in2 => \_gnd_net_\,
            in3 => \N__741\,
            lcout => generated_signal_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1488\,
            ce => 'H',
            sr => \N__1453\
        );

    \fsm_shiftRegs_inst1.current_state_3_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__983\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__765\,
            lcout => \fsm_shiftRegs_inst1.current_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1488\,
            ce => 'H',
            sr => \N__1453\
        );

    \RST_N_ibuf_RNIBJGC_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1268\,
            lcout => \RST_N_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counter_RNO_0_2_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100001000"
        )
    port map (
            in0 => \N__856\,
            in1 => \N__836\,
            in2 => \N__1011\,
            in3 => \N__814\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counter_2_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__717\,
            in3 => \N__1040\,
            lcout => \fsm_shiftRegs_inst1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1495\,
            ce => 'H',
            sr => \N__1456\
        );

    \fsm_shiftRegs_inst1.counter_0_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000001010000"
        )
    port map (
            in0 => \N__857\,
            in1 => \_gnd_net_\,
            in2 => \N__1047\,
            in3 => \N__1008\,
            lcout => \fsm_shiftRegs_inst1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1495\,
            ce => 'H',
            sr => \N__1456\
        );

    \fsm_shiftRegs_inst1.counter_RNIC589_1_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__834\,
            in1 => \N__854\,
            in2 => \_gnd_net_\,
            in3 => \N__1001\,
            lcout => \fsm_shiftRegs_inst1.N_125_1\,
            ltout => \fsm_shiftRegs_inst1.N_125_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_1_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011001110"
        )
    port map (
            in0 => \N__1045\,
            in1 => \N__1224\,
            in2 => \N__864\,
            in3 => \N__815\,
            lcout => \fsm_shiftRegs_inst1.current_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1495\,
            ce => 'H',
            sr => \N__1456\
        );

    \fsm_shiftRegs_inst1.counter_1_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001110000000000"
        )
    port map (
            in0 => \N__1009\,
            in1 => \N__837\,
            in2 => \N__861\,
            in3 => \N__1044\,
            lcout => \fsm_shiftRegs_inst1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1495\,
            ce => 'H',
            sr => \N__1456\
        );

    \fsm_shiftRegs_inst1.counter_RNO_0_3_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__855\,
            in1 => \N__835\,
            in2 => \N__1010\,
            in3 => \N__813\,
            lcout => \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counterDYN_RNO_0_3_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__950\,
            in1 => \N__922\,
            in2 => \N__780\,
            in3 => \N__976\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counterDYN_3_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__798\,
            in3 => \N__1331\,
            lcout => \fsm_shiftRegs_inst1.counterDYNZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1493\,
            ce => 'H',
            sr => \N__1454\
        );

    \fsm_shiftRegs_inst1.counterDYN_0_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__1329\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__980\,
            lcout => \fsm_shiftRegs_inst1.counterDYNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1493\,
            ce => 'H',
            sr => \N__1454\
        );

    \fsm_shiftRegs_inst1.current_state_RNO_0_2_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__923\,
            in1 => \N__951\,
            in2 => \N__984\,
            in3 => \N__779\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_2_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__1330\,
            in1 => \N__795\,
            in2 => \N__789\,
            in3 => \N__786\,
            lcout => \fsm_shiftRegs_inst1.current_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1493\,
            ce => 'H',
            sr => \N__1454\
        );

    \fsm_shiftRegs_inst1.current_state_RNO_0_3_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__921\,
            in1 => \N__1328\,
            in2 => \N__954\,
            in3 => \N__775\,
            lcout => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counterDYN_2_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100100011000000"
        )
    port map (
            in0 => \N__952\,
            in1 => \N__1334\,
            in2 => \N__927\,
            in3 => \N__981\,
            lcout => \fsm_shiftRegs_inst1.counterDYNZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1493\,
            ce => 'H',
            sr => \N__1454\
        );

    \fsm_shiftRegs_inst1.bit_sequence_15_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1212\,
            in2 => \_gnd_net_\,
            in3 => \N__900\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1491\,
            ce => \N__1286\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_14_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__1215\,
            in1 => \N__894\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1491\,
            ce => \N__1286\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_13_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1211\,
            in2 => \_gnd_net_\,
            in3 => \N__888\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1491\,
            ce => \N__1286\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_12_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__1214\,
            in1 => \N__882\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1491\,
            ce => \N__1286\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_11_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1210\,
            in2 => \_gnd_net_\,
            in3 => \N__876\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1491\,
            ce => \N__1286\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_10_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__1213\,
            in1 => \N__1065\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1491\,
            ce => \N__1286\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_6_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__1217\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__870\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1489\,
            ce => \N__1287\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_5_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1083\,
            in2 => \_gnd_net_\,
            in3 => \N__1220\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1489\,
            ce => \N__1287\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_7_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__1218\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1095\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1489\,
            ce => \N__1287\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_3_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1154\,
            in2 => \_gnd_net_\,
            in3 => \N__1219\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1489\,
            ce => \N__1287\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_4_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__1216\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1089\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1489\,
            ce => \N__1287\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_8_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1077\,
            in2 => \_gnd_net_\,
            in3 => \N__1221\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1489\,
            ce => \N__1287\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_9_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1071\,
            in2 => \_gnd_net_\,
            in3 => \N__1222\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1489\,
            ce => \N__1287\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.en_fin_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__1430\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ENFIN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1487\,
            ce => 'H',
            sr => \N__1452\
        );

    \fsm_shiftRegs_inst1.counter_3_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1046\,
            in2 => \_gnd_net_\,
            in3 => \N__1017\,
            lcout => \fsm_shiftRegs_inst1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1496\,
            ce => 'H',
            sr => \N__1457\
        );

    \fsm_shiftRegs_inst1.counterDYN_1_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__1332\,
            in1 => \N__982\,
            in2 => \_gnd_net_\,
            in3 => \N__953\,
            lcout => \fsm_shiftRegs_inst1.counterDYNZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1496\,
            ce => 'H',
            sr => \N__1457\
        );

    \fsm_shiftRegs_inst1.current_state_RNO_0_4_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__1116\,
            in1 => \N__1133\,
            in2 => \N__1605\,
            in3 => \N__1568\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_4_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111011101110"
        )
    port map (
            in0 => \N__1428\,
            in1 => \N__1365\,
            in2 => \N__1350\,
            in3 => \N__1344\,
            lcout => \fsm_shiftRegs_inst1.current_stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1494\,
            ce => 'H',
            sr => \N__1455\
        );

    \fsm_shiftRegs_inst1.current_state_RNO_0_0_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__1601\,
            in1 => \N__1112\,
            in2 => \_gnd_net_\,
            in3 => \N__1567\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_0_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__1134\,
            in1 => \N__1429\,
            in2 => \N__1347\,
            in3 => \N__1343\,
            lcout => \fsm_shiftRegs_inst1.current_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1494\,
            ce => 'H',
            sr => \N__1455\
        );

    \fsm_shiftRegs_inst1.counter2_RNITAO81_7_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1508\,
            in1 => \N__1583\,
            in2 => \N__1548\,
            in3 => \N__1526\,
            lcout => \fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_RNO_0_2_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__1326\,
            in1 => \N__1205\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_shiftRegs_inst1.N_122_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_RNI333L_2_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__1206\,
            in1 => \N__1327\,
            in2 => \_gnd_net_\,
            in3 => \N__1263\,
            lcout => \fsm_shiftRegs_inst1.un1_current_state4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_2_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__1269\,
            in1 => \N__1155\,
            in2 => \_gnd_net_\,
            in3 => \N__1223\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1492\,
            ce => \N__1143\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counter2_0_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1392\,
            in1 => \N__1132\,
            in2 => \_gnd_net_\,
            in3 => \N__1119\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_11_0_\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_0\,
            clk => \N__1497\,
            ce => 'H',
            sr => \N__1458\
        );

    \fsm_shiftRegs_inst1.counter2_1_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1388\,
            in1 => \N__1111\,
            in2 => \_gnd_net_\,
            in3 => \N__1608\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_1\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_0\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_1\,
            clk => \N__1497\,
            ce => 'H',
            sr => \N__1458\
        );

    \fsm_shiftRegs_inst1.counter2_2_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1393\,
            in1 => \N__1600\,
            in2 => \_gnd_net_\,
            in3 => \N__1587\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_2\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_1\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_2\,
            clk => \N__1497\,
            ce => 'H',
            sr => \N__1458\
        );

    \fsm_shiftRegs_inst1.counter2_3_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1389\,
            in1 => \N__1584\,
            in2 => \_gnd_net_\,
            in3 => \N__1572\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_3\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_2\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_3\,
            clk => \N__1497\,
            ce => 'H',
            sr => \N__1458\
        );

    \fsm_shiftRegs_inst1.counter2_4_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__1394\,
            in1 => \_gnd_net_\,
            in2 => \N__1569\,
            in3 => \N__1551\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_4\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_3\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_4\,
            clk => \N__1497\,
            ce => 'H',
            sr => \N__1458\
        );

    \fsm_shiftRegs_inst1.counter2_5_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1390\,
            in1 => \N__1547\,
            in2 => \_gnd_net_\,
            in3 => \N__1533\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_5\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_4\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_5\,
            clk => \N__1497\,
            ce => 'H',
            sr => \N__1458\
        );

    \fsm_shiftRegs_inst1.counter2_6_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__1395\,
            in1 => \_gnd_net_\,
            in2 => \N__1530\,
            in3 => \N__1515\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_6\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_5\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_6\,
            clk => \N__1497\,
            ce => 'H',
            sr => \N__1458\
        );

    \fsm_shiftRegs_inst1.counter2_7_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1391\,
            in1 => \N__1509\,
            in2 => \_gnd_net_\,
            in3 => \N__1512\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1497\,
            ce => 'H',
            sr => \N__1458\
        );

    \fsm_shiftRegs_inst1.current_state_RNIVA94_4_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1421\,
            lcout => \fsm_shiftRegs_inst1.current_state_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
