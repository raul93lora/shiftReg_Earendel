-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 19 2025 11:24:18

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    SDO_signal_out : out std_logic;
    RST_N : in std_logic;
    CLK_uC : in std_logic;
    CLK : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__6294\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3507\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3333\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3303\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3219\ : std_logic;
signal \N__3216\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3144\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \RST_N_c\ : std_logic;
signal \RST_N_c_i\ : std_logic;
signal \fsm_ctrl_inst1.current_state_i_0\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_58\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_57\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_6\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_84\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_85\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_86\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_1\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_2\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_5\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_3\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_4\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_56\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_59\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_55\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_7\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_8\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_9\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_10\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_83\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_42\ : std_logic;
signal \bfn_3_20_0_\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_cry_0\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_cry_1\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_cry_2\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_cry_3\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_9\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_6\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_7\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_8\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_12\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_10\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_11\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_13\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_14\ : std_logic;
signal \fsm_ctrl_inst1.current_state_i_1\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_75\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_76\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_77\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_11\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_54\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_60\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_61\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_78\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_79\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_80\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_4\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_5\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_53\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_37\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_81\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_82\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_3\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_1\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_2\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_38\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_39\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_40\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_41\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_43\ : std_logic;
signal \fsm_ctrl_inst1.g0_0_2_0_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_s_3\ : std_logic;
signal \fsm_ctrl_inst1.g0_0_2_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_s_4\ : std_logic;
signal \fsm_ctrl_inst1.g0_0_3_1\ : std_logic;
signal \fsm_ctrl_inst1.g0_0_2_1\ : std_logic;
signal \fsm_ctrl_inst1.current_state_20_d_i_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_s_2\ : std_logic;
signal \fsm_ctrl_inst1.N_93_0_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.counter_idlee_0_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_s_1\ : std_logic;
signal \fsm_ctrl_inst1.g0_0_3_2\ : std_logic;
signal \fsm_ctrl_inst1.g0_0_2_2\ : std_logic;
signal \fsm_ctrl_inst1.current_state_20_d_i\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_15\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_87\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_67\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_64\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_65\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_66\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_68\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_69\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_70\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_73\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_74\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_71\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_72\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_18\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_17\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_16\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_14\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_15\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_62\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_63\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_21\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_22\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_48\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_26\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_12\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_13\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_49\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_50\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_47\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_25\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_44\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_51\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_52\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_23\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_24\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_45\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_46\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_27\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_28\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_33\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_29\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_34\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_30\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_35\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_36\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_31\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_32\ : std_logic;
signal \fsm_ctrl_inst1.counter_idleZ0Z_1\ : std_logic;
signal \fsm_ctrl_inst1.counter_idleZ0Z_3\ : std_logic;
signal \fsm_ctrl_inst1.counter_idleZ0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.current_state_RNO_2Z0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.g0_0_3_0\ : std_logic;
signal \fsm_ctrl_inst1.counter_idleZ1Z_4\ : std_logic;
signal \fsm_ctrl_inst1.counter_idleZ0Z_2\ : std_logic;
signal \fsm_ctrl_inst1.g0_0_3\ : std_logic;
signal \fsm_ctrl_inst1.counter_din_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.current_state_RNO_3Z0Z_0_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.current_state_RNO_1Z0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.counter_dinZ0Z_2\ : std_logic;
signal \fsm_ctrl_inst1.counter_dinZ0Z_3\ : std_logic;
signal \fsm_ctrl_inst1.counter_dinZ0Z_1\ : std_logic;
signal \fsm_ctrl_inst1.counter_dinZ0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.o2_cascade_\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_19\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_20\ : std_logic;
signal \fsm_ctrl_inst1.current_state_i_g_0\ : std_logic;
signal \SDO_signal_out_c\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_14\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_15\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_12\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_13\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_10\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_11\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSR_cnv_x0Z0Z_0_cascade_\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSR_cnv_x1Z0Z_0\ : std_logic;
signal \CLK_uC_c\ : std_logic;
signal \fsm_ctrl_inst1_SCLK_i\ : std_logic;
signal fsm_ctrl_inst1_current_state_1 : std_logic;
signal \config_register_latched_dec_inst1.STATSR_cnv_x1Z0Z_0_cascade_\ : std_logic;
signal \config_register_latched_dec_inst1.STATSR_cnv_x0Z0Z_0\ : std_logic;
signal \STATSR_cnv_ns_0\ : std_logic;
signal fsm_ctrl_inst1_current_state_0 : std_logic;
signal \SEL_REG\ : std_logic;
signal \MOSI\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_0\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_1\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_2\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_3\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_1\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_2\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_3\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_87\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_9\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_6\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_7\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_8\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_4\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_5\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSR_cnv_nsZ0Z_0\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_4\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_5\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_86\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_6\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_7\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_8\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_84\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_85\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_9\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_10\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_11\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_83\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_12\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_81\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_82\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_13\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_80\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_79\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_77\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_78\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_14\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_75\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_76\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_74\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_15\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_16\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_73\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_17\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_18\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_71\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_72\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_70\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_68\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_69\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_67\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_66\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_19\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_20\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_41\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_40\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_42\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_43\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_44\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_45\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_21\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_65\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_36\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_35\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_37\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_38\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_39\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_46\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_47\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_22\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_48\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_23\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_49\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_52\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_50\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_51\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_64\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_63\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_53\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_61\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_62\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_30\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_34\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_31\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_32\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_33\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_26\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_24\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_25\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_27\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_28\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_29\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_60\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_54\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_59\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_57\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_58\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_55\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_56\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \CLK_0_c_g\ : std_logic;
signal \N_218_g\ : std_logic;
signal \RST_N_c_i_g\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \CLK_uC_wire\ : std_logic;
signal \RST_N_wire\ : std_logic;
signal \SDO_signal_out_wire\ : std_logic;

begin
    \CLK_wire\ <= CLK;
    \CLK_uC_wire\ <= CLK_uC;
    \RST_N_wire\ <= RST_N;
    SDO_signal_out <= \SDO_signal_out_wire\;

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6292\,
            GLOBALBUFFEROUTPUT => \CLK_0_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6294\,
            DIN => \N__6293\,
            DOUT => \N__6292\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6294\,
            PADOUT => \N__6293\,
            PADIN => \N__6292\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_uC_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6283\,
            DIN => \N__6282\,
            DOUT => \N__6281\,
            PACKAGEPIN => \CLK_uC_wire\
        );

    \CLK_uC_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6283\,
            PADOUT => \N__6282\,
            PADIN => \N__6281\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK_uC_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RST_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6274\,
            DIN => \N__6273\,
            DOUT => \N__6272\,
            PACKAGEPIN => \RST_N_wire\
        );

    \RST_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6274\,
            PADOUT => \N__6273\,
            PADIN => \N__6272\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RST_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SDO_signal_out_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6265\,
            DIN => \N__6264\,
            DOUT => \N__6263\,
            PACKAGEPIN => \SDO_signal_out_wire\
        );

    \SDO_signal_out_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6265\,
            PADOUT => \N__6264\,
            PADIN => \N__6263\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4149\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1304\ : InMux
    port map (
            O => \N__6246\,
            I => \N__6243\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__6243\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_27\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6240\,
            I => \N__6237\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__6237\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_28\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6234\,
            I => \N__6231\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6231\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_29\
        );

    \I__1298\ : InMux
    port map (
            O => \N__6228\,
            I => \N__6225\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__6225\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_60\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6222\,
            I => \N__6219\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__6219\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_54\
        );

    \I__1294\ : InMux
    port map (
            O => \N__6216\,
            I => \N__6213\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6213\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_59\
        );

    \I__1292\ : InMux
    port map (
            O => \N__6210\,
            I => \N__6207\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__6207\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_57\
        );

    \I__1290\ : InMux
    port map (
            O => \N__6204\,
            I => \N__6201\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__6201\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_58\
        );

    \I__1288\ : InMux
    port map (
            O => \N__6198\,
            I => \N__6195\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__6195\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_55\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6192\,
            I => \N__6189\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__6189\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_56\
        );

    \I__1284\ : ClkMux
    port map (
            O => \N__6186\,
            I => \N__5982\
        );

    \I__1283\ : ClkMux
    port map (
            O => \N__6185\,
            I => \N__5982\
        );

    \I__1282\ : ClkMux
    port map (
            O => \N__6184\,
            I => \N__5982\
        );

    \I__1281\ : ClkMux
    port map (
            O => \N__6183\,
            I => \N__5982\
        );

    \I__1280\ : ClkMux
    port map (
            O => \N__6182\,
            I => \N__5982\
        );

    \I__1279\ : ClkMux
    port map (
            O => \N__6181\,
            I => \N__5982\
        );

    \I__1278\ : ClkMux
    port map (
            O => \N__6180\,
            I => \N__5982\
        );

    \I__1277\ : ClkMux
    port map (
            O => \N__6179\,
            I => \N__5982\
        );

    \I__1276\ : ClkMux
    port map (
            O => \N__6178\,
            I => \N__5982\
        );

    \I__1275\ : ClkMux
    port map (
            O => \N__6177\,
            I => \N__5982\
        );

    \I__1274\ : ClkMux
    port map (
            O => \N__6176\,
            I => \N__5982\
        );

    \I__1273\ : ClkMux
    port map (
            O => \N__6175\,
            I => \N__5982\
        );

    \I__1272\ : ClkMux
    port map (
            O => \N__6174\,
            I => \N__5982\
        );

    \I__1271\ : ClkMux
    port map (
            O => \N__6173\,
            I => \N__5982\
        );

    \I__1270\ : ClkMux
    port map (
            O => \N__6172\,
            I => \N__5982\
        );

    \I__1269\ : ClkMux
    port map (
            O => \N__6171\,
            I => \N__5982\
        );

    \I__1268\ : ClkMux
    port map (
            O => \N__6170\,
            I => \N__5982\
        );

    \I__1267\ : ClkMux
    port map (
            O => \N__6169\,
            I => \N__5982\
        );

    \I__1266\ : ClkMux
    port map (
            O => \N__6168\,
            I => \N__5982\
        );

    \I__1265\ : ClkMux
    port map (
            O => \N__6167\,
            I => \N__5982\
        );

    \I__1264\ : ClkMux
    port map (
            O => \N__6166\,
            I => \N__5982\
        );

    \I__1263\ : ClkMux
    port map (
            O => \N__6165\,
            I => \N__5982\
        );

    \I__1262\ : ClkMux
    port map (
            O => \N__6164\,
            I => \N__5982\
        );

    \I__1261\ : ClkMux
    port map (
            O => \N__6163\,
            I => \N__5982\
        );

    \I__1260\ : ClkMux
    port map (
            O => \N__6162\,
            I => \N__5982\
        );

    \I__1259\ : ClkMux
    port map (
            O => \N__6161\,
            I => \N__5982\
        );

    \I__1258\ : ClkMux
    port map (
            O => \N__6160\,
            I => \N__5982\
        );

    \I__1257\ : ClkMux
    port map (
            O => \N__6159\,
            I => \N__5982\
        );

    \I__1256\ : ClkMux
    port map (
            O => \N__6158\,
            I => \N__5982\
        );

    \I__1255\ : ClkMux
    port map (
            O => \N__6157\,
            I => \N__5982\
        );

    \I__1254\ : ClkMux
    port map (
            O => \N__6156\,
            I => \N__5982\
        );

    \I__1253\ : ClkMux
    port map (
            O => \N__6155\,
            I => \N__5982\
        );

    \I__1252\ : ClkMux
    port map (
            O => \N__6154\,
            I => \N__5982\
        );

    \I__1251\ : ClkMux
    port map (
            O => \N__6153\,
            I => \N__5982\
        );

    \I__1250\ : ClkMux
    port map (
            O => \N__6152\,
            I => \N__5982\
        );

    \I__1249\ : ClkMux
    port map (
            O => \N__6151\,
            I => \N__5982\
        );

    \I__1248\ : ClkMux
    port map (
            O => \N__6150\,
            I => \N__5982\
        );

    \I__1247\ : ClkMux
    port map (
            O => \N__6149\,
            I => \N__5982\
        );

    \I__1246\ : ClkMux
    port map (
            O => \N__6148\,
            I => \N__5982\
        );

    \I__1245\ : ClkMux
    port map (
            O => \N__6147\,
            I => \N__5982\
        );

    \I__1244\ : ClkMux
    port map (
            O => \N__6146\,
            I => \N__5982\
        );

    \I__1243\ : ClkMux
    port map (
            O => \N__6145\,
            I => \N__5982\
        );

    \I__1242\ : ClkMux
    port map (
            O => \N__6144\,
            I => \N__5982\
        );

    \I__1241\ : ClkMux
    port map (
            O => \N__6143\,
            I => \N__5982\
        );

    \I__1240\ : ClkMux
    port map (
            O => \N__6142\,
            I => \N__5982\
        );

    \I__1239\ : ClkMux
    port map (
            O => \N__6141\,
            I => \N__5982\
        );

    \I__1238\ : ClkMux
    port map (
            O => \N__6140\,
            I => \N__5982\
        );

    \I__1237\ : ClkMux
    port map (
            O => \N__6139\,
            I => \N__5982\
        );

    \I__1236\ : ClkMux
    port map (
            O => \N__6138\,
            I => \N__5982\
        );

    \I__1235\ : ClkMux
    port map (
            O => \N__6137\,
            I => \N__5982\
        );

    \I__1234\ : ClkMux
    port map (
            O => \N__6136\,
            I => \N__5982\
        );

    \I__1233\ : ClkMux
    port map (
            O => \N__6135\,
            I => \N__5982\
        );

    \I__1232\ : ClkMux
    port map (
            O => \N__6134\,
            I => \N__5982\
        );

    \I__1231\ : ClkMux
    port map (
            O => \N__6133\,
            I => \N__5982\
        );

    \I__1230\ : ClkMux
    port map (
            O => \N__6132\,
            I => \N__5982\
        );

    \I__1229\ : ClkMux
    port map (
            O => \N__6131\,
            I => \N__5982\
        );

    \I__1228\ : ClkMux
    port map (
            O => \N__6130\,
            I => \N__5982\
        );

    \I__1227\ : ClkMux
    port map (
            O => \N__6129\,
            I => \N__5982\
        );

    \I__1226\ : ClkMux
    port map (
            O => \N__6128\,
            I => \N__5982\
        );

    \I__1225\ : ClkMux
    port map (
            O => \N__6127\,
            I => \N__5982\
        );

    \I__1224\ : ClkMux
    port map (
            O => \N__6126\,
            I => \N__5982\
        );

    \I__1223\ : ClkMux
    port map (
            O => \N__6125\,
            I => \N__5982\
        );

    \I__1222\ : ClkMux
    port map (
            O => \N__6124\,
            I => \N__5982\
        );

    \I__1221\ : ClkMux
    port map (
            O => \N__6123\,
            I => \N__5982\
        );

    \I__1220\ : ClkMux
    port map (
            O => \N__6122\,
            I => \N__5982\
        );

    \I__1219\ : ClkMux
    port map (
            O => \N__6121\,
            I => \N__5982\
        );

    \I__1218\ : ClkMux
    port map (
            O => \N__6120\,
            I => \N__5982\
        );

    \I__1217\ : ClkMux
    port map (
            O => \N__6119\,
            I => \N__5982\
        );

    \I__1216\ : GlobalMux
    port map (
            O => \N__5982\,
            I => \N__5979\
        );

    \I__1215\ : gio2CtrlBuf
    port map (
            O => \N__5979\,
            I => \CLK_0_c_g\
        );

    \I__1214\ : CEMux
    port map (
            O => \N__5976\,
            I => \N__5874\
        );

    \I__1213\ : CEMux
    port map (
            O => \N__5975\,
            I => \N__5874\
        );

    \I__1212\ : CEMux
    port map (
            O => \N__5974\,
            I => \N__5874\
        );

    \I__1211\ : CEMux
    port map (
            O => \N__5973\,
            I => \N__5874\
        );

    \I__1210\ : CEMux
    port map (
            O => \N__5972\,
            I => \N__5874\
        );

    \I__1209\ : CEMux
    port map (
            O => \N__5971\,
            I => \N__5874\
        );

    \I__1208\ : CEMux
    port map (
            O => \N__5970\,
            I => \N__5874\
        );

    \I__1207\ : CEMux
    port map (
            O => \N__5969\,
            I => \N__5874\
        );

    \I__1206\ : CEMux
    port map (
            O => \N__5968\,
            I => \N__5874\
        );

    \I__1205\ : CEMux
    port map (
            O => \N__5967\,
            I => \N__5874\
        );

    \I__1204\ : CEMux
    port map (
            O => \N__5966\,
            I => \N__5874\
        );

    \I__1203\ : CEMux
    port map (
            O => \N__5965\,
            I => \N__5874\
        );

    \I__1202\ : CEMux
    port map (
            O => \N__5964\,
            I => \N__5874\
        );

    \I__1201\ : CEMux
    port map (
            O => \N__5963\,
            I => \N__5874\
        );

    \I__1200\ : CEMux
    port map (
            O => \N__5962\,
            I => \N__5874\
        );

    \I__1199\ : CEMux
    port map (
            O => \N__5961\,
            I => \N__5874\
        );

    \I__1198\ : CEMux
    port map (
            O => \N__5960\,
            I => \N__5874\
        );

    \I__1197\ : CEMux
    port map (
            O => \N__5959\,
            I => \N__5874\
        );

    \I__1196\ : CEMux
    port map (
            O => \N__5958\,
            I => \N__5874\
        );

    \I__1195\ : CEMux
    port map (
            O => \N__5957\,
            I => \N__5874\
        );

    \I__1194\ : CEMux
    port map (
            O => \N__5956\,
            I => \N__5874\
        );

    \I__1193\ : CEMux
    port map (
            O => \N__5955\,
            I => \N__5874\
        );

    \I__1192\ : CEMux
    port map (
            O => \N__5954\,
            I => \N__5874\
        );

    \I__1191\ : CEMux
    port map (
            O => \N__5953\,
            I => \N__5874\
        );

    \I__1190\ : CEMux
    port map (
            O => \N__5952\,
            I => \N__5874\
        );

    \I__1189\ : CEMux
    port map (
            O => \N__5951\,
            I => \N__5874\
        );

    \I__1188\ : CEMux
    port map (
            O => \N__5950\,
            I => \N__5874\
        );

    \I__1187\ : CEMux
    port map (
            O => \N__5949\,
            I => \N__5874\
        );

    \I__1186\ : CEMux
    port map (
            O => \N__5948\,
            I => \N__5874\
        );

    \I__1185\ : CEMux
    port map (
            O => \N__5947\,
            I => \N__5874\
        );

    \I__1184\ : CEMux
    port map (
            O => \N__5946\,
            I => \N__5874\
        );

    \I__1183\ : CEMux
    port map (
            O => \N__5945\,
            I => \N__5874\
        );

    \I__1182\ : CEMux
    port map (
            O => \N__5944\,
            I => \N__5874\
        );

    \I__1181\ : CEMux
    port map (
            O => \N__5943\,
            I => \N__5874\
        );

    \I__1180\ : GlobalMux
    port map (
            O => \N__5874\,
            I => \N__5871\
        );

    \I__1179\ : gio2CtrlBuf
    port map (
            O => \N__5871\,
            I => \N_218_g\
        );

    \I__1178\ : SRMux
    port map (
            O => \N__5868\,
            I => \N__5664\
        );

    \I__1177\ : SRMux
    port map (
            O => \N__5867\,
            I => \N__5664\
        );

    \I__1176\ : SRMux
    port map (
            O => \N__5866\,
            I => \N__5664\
        );

    \I__1175\ : SRMux
    port map (
            O => \N__5865\,
            I => \N__5664\
        );

    \I__1174\ : SRMux
    port map (
            O => \N__5864\,
            I => \N__5664\
        );

    \I__1173\ : SRMux
    port map (
            O => \N__5863\,
            I => \N__5664\
        );

    \I__1172\ : SRMux
    port map (
            O => \N__5862\,
            I => \N__5664\
        );

    \I__1171\ : SRMux
    port map (
            O => \N__5861\,
            I => \N__5664\
        );

    \I__1170\ : SRMux
    port map (
            O => \N__5860\,
            I => \N__5664\
        );

    \I__1169\ : SRMux
    port map (
            O => \N__5859\,
            I => \N__5664\
        );

    \I__1168\ : SRMux
    port map (
            O => \N__5858\,
            I => \N__5664\
        );

    \I__1167\ : SRMux
    port map (
            O => \N__5857\,
            I => \N__5664\
        );

    \I__1166\ : SRMux
    port map (
            O => \N__5856\,
            I => \N__5664\
        );

    \I__1165\ : SRMux
    port map (
            O => \N__5855\,
            I => \N__5664\
        );

    \I__1164\ : SRMux
    port map (
            O => \N__5854\,
            I => \N__5664\
        );

    \I__1163\ : SRMux
    port map (
            O => \N__5853\,
            I => \N__5664\
        );

    \I__1162\ : SRMux
    port map (
            O => \N__5852\,
            I => \N__5664\
        );

    \I__1161\ : SRMux
    port map (
            O => \N__5851\,
            I => \N__5664\
        );

    \I__1160\ : SRMux
    port map (
            O => \N__5850\,
            I => \N__5664\
        );

    \I__1159\ : SRMux
    port map (
            O => \N__5849\,
            I => \N__5664\
        );

    \I__1158\ : SRMux
    port map (
            O => \N__5848\,
            I => \N__5664\
        );

    \I__1157\ : SRMux
    port map (
            O => \N__5847\,
            I => \N__5664\
        );

    \I__1156\ : SRMux
    port map (
            O => \N__5846\,
            I => \N__5664\
        );

    \I__1155\ : SRMux
    port map (
            O => \N__5845\,
            I => \N__5664\
        );

    \I__1154\ : SRMux
    port map (
            O => \N__5844\,
            I => \N__5664\
        );

    \I__1153\ : SRMux
    port map (
            O => \N__5843\,
            I => \N__5664\
        );

    \I__1152\ : SRMux
    port map (
            O => \N__5842\,
            I => \N__5664\
        );

    \I__1151\ : SRMux
    port map (
            O => \N__5841\,
            I => \N__5664\
        );

    \I__1150\ : SRMux
    port map (
            O => \N__5840\,
            I => \N__5664\
        );

    \I__1149\ : SRMux
    port map (
            O => \N__5839\,
            I => \N__5664\
        );

    \I__1148\ : SRMux
    port map (
            O => \N__5838\,
            I => \N__5664\
        );

    \I__1147\ : SRMux
    port map (
            O => \N__5837\,
            I => \N__5664\
        );

    \I__1146\ : SRMux
    port map (
            O => \N__5836\,
            I => \N__5664\
        );

    \I__1145\ : SRMux
    port map (
            O => \N__5835\,
            I => \N__5664\
        );

    \I__1144\ : SRMux
    port map (
            O => \N__5834\,
            I => \N__5664\
        );

    \I__1143\ : SRMux
    port map (
            O => \N__5833\,
            I => \N__5664\
        );

    \I__1142\ : SRMux
    port map (
            O => \N__5832\,
            I => \N__5664\
        );

    \I__1141\ : SRMux
    port map (
            O => \N__5831\,
            I => \N__5664\
        );

    \I__1140\ : SRMux
    port map (
            O => \N__5830\,
            I => \N__5664\
        );

    \I__1139\ : SRMux
    port map (
            O => \N__5829\,
            I => \N__5664\
        );

    \I__1138\ : SRMux
    port map (
            O => \N__5828\,
            I => \N__5664\
        );

    \I__1137\ : SRMux
    port map (
            O => \N__5827\,
            I => \N__5664\
        );

    \I__1136\ : SRMux
    port map (
            O => \N__5826\,
            I => \N__5664\
        );

    \I__1135\ : SRMux
    port map (
            O => \N__5825\,
            I => \N__5664\
        );

    \I__1134\ : SRMux
    port map (
            O => \N__5824\,
            I => \N__5664\
        );

    \I__1133\ : SRMux
    port map (
            O => \N__5823\,
            I => \N__5664\
        );

    \I__1132\ : SRMux
    port map (
            O => \N__5822\,
            I => \N__5664\
        );

    \I__1131\ : SRMux
    port map (
            O => \N__5821\,
            I => \N__5664\
        );

    \I__1130\ : SRMux
    port map (
            O => \N__5820\,
            I => \N__5664\
        );

    \I__1129\ : SRMux
    port map (
            O => \N__5819\,
            I => \N__5664\
        );

    \I__1128\ : SRMux
    port map (
            O => \N__5818\,
            I => \N__5664\
        );

    \I__1127\ : SRMux
    port map (
            O => \N__5817\,
            I => \N__5664\
        );

    \I__1126\ : SRMux
    port map (
            O => \N__5816\,
            I => \N__5664\
        );

    \I__1125\ : SRMux
    port map (
            O => \N__5815\,
            I => \N__5664\
        );

    \I__1124\ : SRMux
    port map (
            O => \N__5814\,
            I => \N__5664\
        );

    \I__1123\ : SRMux
    port map (
            O => \N__5813\,
            I => \N__5664\
        );

    \I__1122\ : SRMux
    port map (
            O => \N__5812\,
            I => \N__5664\
        );

    \I__1121\ : SRMux
    port map (
            O => \N__5811\,
            I => \N__5664\
        );

    \I__1120\ : SRMux
    port map (
            O => \N__5810\,
            I => \N__5664\
        );

    \I__1119\ : SRMux
    port map (
            O => \N__5809\,
            I => \N__5664\
        );

    \I__1118\ : SRMux
    port map (
            O => \N__5808\,
            I => \N__5664\
        );

    \I__1117\ : SRMux
    port map (
            O => \N__5807\,
            I => \N__5664\
        );

    \I__1116\ : SRMux
    port map (
            O => \N__5806\,
            I => \N__5664\
        );

    \I__1115\ : SRMux
    port map (
            O => \N__5805\,
            I => \N__5664\
        );

    \I__1114\ : SRMux
    port map (
            O => \N__5804\,
            I => \N__5664\
        );

    \I__1113\ : SRMux
    port map (
            O => \N__5803\,
            I => \N__5664\
        );

    \I__1112\ : SRMux
    port map (
            O => \N__5802\,
            I => \N__5664\
        );

    \I__1111\ : SRMux
    port map (
            O => \N__5801\,
            I => \N__5664\
        );

    \I__1110\ : GlobalMux
    port map (
            O => \N__5664\,
            I => \N__5661\
        );

    \I__1109\ : gio2CtrlBuf
    port map (
            O => \N__5661\,
            I => \RST_N_c_i_g\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5658\,
            I => \N__5655\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__5655\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_61\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5652\,
            I => \N__5649\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5649\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_62\
        );

    \I__1104\ : InMux
    port map (
            O => \N__5646\,
            I => \N__5643\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5643\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_30\
        );

    \I__1102\ : InMux
    port map (
            O => \N__5640\,
            I => \N__5637\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__5637\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_34\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5634\,
            I => \N__5631\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5631\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_31\
        );

    \I__1098\ : InMux
    port map (
            O => \N__5628\,
            I => \N__5625\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5625\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_32\
        );

    \I__1096\ : InMux
    port map (
            O => \N__5622\,
            I => \N__5619\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__5619\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_33\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5616\,
            I => \N__5613\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__5613\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_26\
        );

    \I__1092\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5607\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5607\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_24\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5604\,
            I => \N__5601\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__5601\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_25\
        );

    \I__1088\ : InMux
    port map (
            O => \N__5598\,
            I => \N__5595\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__5595\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_23\
        );

    \I__1086\ : InMux
    port map (
            O => \N__5592\,
            I => \N__5589\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__5589\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_49\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5586\,
            I => \N__5583\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__5583\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_52\
        );

    \I__1082\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5577\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__5577\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_50\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5574\,
            I => \N__5571\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__5571\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_51\
        );

    \I__1078\ : InMux
    port map (
            O => \N__5568\,
            I => \N__5565\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5565\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_64\
        );

    \I__1076\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5559\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__5559\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_63\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5556\,
            I => \N__5553\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__5553\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_53\
        );

    \I__1072\ : InMux
    port map (
            O => \N__5550\,
            I => \N__5547\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__5547\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_36\
        );

    \I__1070\ : InMux
    port map (
            O => \N__5544\,
            I => \N__5541\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__5541\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_35\
        );

    \I__1068\ : InMux
    port map (
            O => \N__5538\,
            I => \N__5535\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__5535\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_37\
        );

    \I__1066\ : InMux
    port map (
            O => \N__5532\,
            I => \N__5529\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__5529\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_38\
        );

    \I__1064\ : InMux
    port map (
            O => \N__5526\,
            I => \N__5523\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__5523\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_39\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5517\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5517\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_46\
        );

    \I__1060\ : InMux
    port map (
            O => \N__5514\,
            I => \N__5511\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5511\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_47\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5508\,
            I => \N__5505\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__5505\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_22\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5502\,
            I => \N__5499\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__5499\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_48\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5496\,
            I => \N__5493\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__5493\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_19\
        );

    \I__1052\ : InMux
    port map (
            O => \N__5490\,
            I => \N__5487\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__5487\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_20\
        );

    \I__1050\ : InMux
    port map (
            O => \N__5484\,
            I => \N__5481\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__5481\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_41\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5478\,
            I => \N__5475\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__5475\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_40\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5472\,
            I => \N__5469\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__5469\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_42\
        );

    \I__1044\ : InMux
    port map (
            O => \N__5466\,
            I => \N__5463\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__5463\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_43\
        );

    \I__1042\ : InMux
    port map (
            O => \N__5460\,
            I => \N__5457\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__5457\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_44\
        );

    \I__1040\ : InMux
    port map (
            O => \N__5454\,
            I => \N__5451\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__5451\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_45\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5448\,
            I => \N__5445\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__5445\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_21\
        );

    \I__1036\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5439\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__5439\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_65\
        );

    \I__1034\ : InMux
    port map (
            O => \N__5436\,
            I => \N__5433\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__5433\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_18\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5430\,
            I => \N__5427\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__5427\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_71\
        );

    \I__1030\ : InMux
    port map (
            O => \N__5424\,
            I => \N__5421\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__5421\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_72\
        );

    \I__1028\ : InMux
    port map (
            O => \N__5418\,
            I => \N__5415\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__5415\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_70\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5412\,
            I => \N__5409\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__5409\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_68\
        );

    \I__1024\ : InMux
    port map (
            O => \N__5406\,
            I => \N__5403\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__5403\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_69\
        );

    \I__1022\ : InMux
    port map (
            O => \N__5400\,
            I => \N__5397\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__5397\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_67\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5394\,
            I => \N__5391\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__5391\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_66\
        );

    \I__1018\ : InMux
    port map (
            O => \N__5388\,
            I => \N__5385\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__5385\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_77\
        );

    \I__1016\ : InMux
    port map (
            O => \N__5382\,
            I => \N__5379\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5379\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_78\
        );

    \I__1014\ : InMux
    port map (
            O => \N__5376\,
            I => \N__5373\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__5373\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_14\
        );

    \I__1012\ : InMux
    port map (
            O => \N__5370\,
            I => \N__5367\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__5367\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_75\
        );

    \I__1010\ : InMux
    port map (
            O => \N__5364\,
            I => \N__5361\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__5361\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_76\
        );

    \I__1008\ : InMux
    port map (
            O => \N__5358\,
            I => \N__5355\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__5355\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_74\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5352\,
            I => \N__5349\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__5349\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_15\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5346\,
            I => \N__5343\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5343\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_16\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5340\,
            I => \N__5337\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__5337\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_73\
        );

    \I__1000\ : InMux
    port map (
            O => \N__5334\,
            I => \N__5331\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__5331\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_17\
        );

    \I__998\ : InMux
    port map (
            O => \N__5328\,
            I => \N__5325\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__5325\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_10\
        );

    \I__996\ : InMux
    port map (
            O => \N__5322\,
            I => \N__5319\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__5319\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_11\
        );

    \I__994\ : InMux
    port map (
            O => \N__5316\,
            I => \N__5313\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__5313\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_83\
        );

    \I__992\ : InMux
    port map (
            O => \N__5310\,
            I => \N__5307\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__5307\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_12\
        );

    \I__990\ : InMux
    port map (
            O => \N__5304\,
            I => \N__5301\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__5301\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_81\
        );

    \I__988\ : InMux
    port map (
            O => \N__5298\,
            I => \N__5295\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__5295\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_82\
        );

    \I__986\ : InMux
    port map (
            O => \N__5292\,
            I => \N__5289\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__5289\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_13\
        );

    \I__984\ : InMux
    port map (
            O => \N__5286\,
            I => \N__5283\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5283\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_80\
        );

    \I__982\ : InMux
    port map (
            O => \N__5280\,
            I => \N__5277\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5277\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_79\
        );

    \I__980\ : InMux
    port map (
            O => \N__5274\,
            I => \N__5271\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__5271\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_4\
        );

    \I__978\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5265\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__5265\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_5\
        );

    \I__976\ : InMux
    port map (
            O => \N__5262\,
            I => \N__5259\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__5259\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_86\
        );

    \I__974\ : InMux
    port map (
            O => \N__5256\,
            I => \N__5253\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__5253\,
            I => \N__5250\
        );

    \I__972\ : Odrv4
    port map (
            O => \N__5250\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_6\
        );

    \I__971\ : InMux
    port map (
            O => \N__5247\,
            I => \N__5244\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__5244\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_7\
        );

    \I__969\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5238\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5238\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_8\
        );

    \I__967\ : InMux
    port map (
            O => \N__5235\,
            I => \N__5232\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5232\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_84\
        );

    \I__965\ : InMux
    port map (
            O => \N__5229\,
            I => \N__5226\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__5226\,
            I => \N__5223\
        );

    \I__963\ : Odrv4
    port map (
            O => \N__5223\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_85\
        );

    \I__962\ : InMux
    port map (
            O => \N__5220\,
            I => \N__5217\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__5217\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_9\
        );

    \I__960\ : InMux
    port map (
            O => \N__5214\,
            I => \N__5211\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__5211\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_2\
        );

    \I__958\ : InMux
    port map (
            O => \N__5208\,
            I => \N__5205\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__5205\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_3\
        );

    \I__956\ : InMux
    port map (
            O => \N__5202\,
            I => \N__5199\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__5199\,
            I => \N__5196\
        );

    \I__954\ : Odrv12
    port map (
            O => \N__5196\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_87\
        );

    \I__953\ : InMux
    port map (
            O => \N__5193\,
            I => \N__5190\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__5190\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_9\
        );

    \I__951\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5184\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__5184\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_6\
        );

    \I__949\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5178\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__5178\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_7\
        );

    \I__947\ : InMux
    port map (
            O => \N__5175\,
            I => \N__5172\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__5172\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_8\
        );

    \I__945\ : InMux
    port map (
            O => \N__5169\,
            I => \N__5166\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__5166\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_4\
        );

    \I__943\ : InMux
    port map (
            O => \N__5163\,
            I => \N__5160\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__5160\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_5\
        );

    \I__941\ : CEMux
    port map (
            O => \N__5157\,
            I => \N__5154\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__5154\,
            I => \N__5149\
        );

    \I__939\ : CEMux
    port map (
            O => \N__5153\,
            I => \N__5146\
        );

    \I__938\ : CEMux
    port map (
            O => \N__5152\,
            I => \N__5142\
        );

    \I__937\ : Span4Mux_h
    port map (
            O => \N__5149\,
            I => \N__5137\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__5146\,
            I => \N__5137\
        );

    \I__935\ : CEMux
    port map (
            O => \N__5145\,
            I => \N__5134\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5142\,
            I => \N__5131\
        );

    \I__933\ : Span4Mux_v
    port map (
            O => \N__5137\,
            I => \N__5126\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__5134\,
            I => \N__5126\
        );

    \I__931\ : Span4Mux_h
    port map (
            O => \N__5131\,
            I => \N__5123\
        );

    \I__930\ : Span4Mux_v
    port map (
            O => \N__5126\,
            I => \N__5120\
        );

    \I__929\ : Odrv4
    port map (
            O => \N__5123\,
            I => \config_register_latched_dec_inst1.DYNSR_cnv_nsZ0Z_0\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__5120\,
            I => \config_register_latched_dec_inst1.DYNSR_cnv_nsZ0Z_0\
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__5115\,
            I => \N__5109\
        );

    \I__926\ : InMux
    port map (
            O => \N__5114\,
            I => \N__5106\
        );

    \I__925\ : InMux
    port map (
            O => \N__5113\,
            I => \N__5099\
        );

    \I__924\ : InMux
    port map (
            O => \N__5112\,
            I => \N__5099\
        );

    \I__923\ : InMux
    port map (
            O => \N__5109\,
            I => \N__5099\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__5106\,
            I => \N__5094\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__5099\,
            I => \N__5094\
        );

    \I__920\ : Span4Mux_v
    port map (
            O => \N__5094\,
            I => \N__5090\
        );

    \I__919\ : InMux
    port map (
            O => \N__5093\,
            I => \N__5087\
        );

    \I__918\ : Span4Mux_h
    port map (
            O => \N__5090\,
            I => \N__5084\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__5087\,
            I => \N__5081\
        );

    \I__916\ : Odrv4
    port map (
            O => \N__5084\,
            I => \CLK_uC_c\
        );

    \I__915\ : Odrv12
    port map (
            O => \N__5081\,
            I => \CLK_uC_c\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__5076\,
            I => \N__5070\
        );

    \I__913\ : InMux
    port map (
            O => \N__5075\,
            I => \N__5063\
        );

    \I__912\ : InMux
    port map (
            O => \N__5074\,
            I => \N__5063\
        );

    \I__911\ : InMux
    port map (
            O => \N__5073\,
            I => \N__5063\
        );

    \I__910\ : InMux
    port map (
            O => \N__5070\,
            I => \N__5060\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5063\,
            I => \fsm_ctrl_inst1_SCLK_i\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__5060\,
            I => \fsm_ctrl_inst1_SCLK_i\
        );

    \I__907\ : InMux
    port map (
            O => \N__5055\,
            I => \N__5040\
        );

    \I__906\ : InMux
    port map (
            O => \N__5054\,
            I => \N__5040\
        );

    \I__905\ : InMux
    port map (
            O => \N__5053\,
            I => \N__5025\
        );

    \I__904\ : InMux
    port map (
            O => \N__5052\,
            I => \N__5025\
        );

    \I__903\ : InMux
    port map (
            O => \N__5051\,
            I => \N__5025\
        );

    \I__902\ : InMux
    port map (
            O => \N__5050\,
            I => \N__5025\
        );

    \I__901\ : InMux
    port map (
            O => \N__5049\,
            I => \N__5025\
        );

    \I__900\ : InMux
    port map (
            O => \N__5048\,
            I => \N__5019\
        );

    \I__899\ : InMux
    port map (
            O => \N__5047\,
            I => \N__5012\
        );

    \I__898\ : InMux
    port map (
            O => \N__5046\,
            I => \N__5012\
        );

    \I__897\ : InMux
    port map (
            O => \N__5045\,
            I => \N__5012\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5040\,
            I => \N__4980\
        );

    \I__895\ : InMux
    port map (
            O => \N__5039\,
            I => \N__4973\
        );

    \I__894\ : InMux
    port map (
            O => \N__5038\,
            I => \N__4973\
        );

    \I__893\ : InMux
    port map (
            O => \N__5037\,
            I => \N__4973\
        );

    \I__892\ : InMux
    port map (
            O => \N__5036\,
            I => \N__4957\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__5025\,
            I => \N__4939\
        );

    \I__890\ : InMux
    port map (
            O => \N__5024\,
            I => \N__4932\
        );

    \I__889\ : InMux
    port map (
            O => \N__5023\,
            I => \N__4932\
        );

    \I__888\ : InMux
    port map (
            O => \N__5022\,
            I => \N__4932\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5019\,
            I => \N__4927\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__5012\,
            I => \N__4927\
        );

    \I__885\ : InMux
    port map (
            O => \N__5011\,
            I => \N__4922\
        );

    \I__884\ : InMux
    port map (
            O => \N__5010\,
            I => \N__4922\
        );

    \I__883\ : InMux
    port map (
            O => \N__5009\,
            I => \N__4911\
        );

    \I__882\ : InMux
    port map (
            O => \N__5008\,
            I => \N__4911\
        );

    \I__881\ : InMux
    port map (
            O => \N__5007\,
            I => \N__4911\
        );

    \I__880\ : InMux
    port map (
            O => \N__5006\,
            I => \N__4911\
        );

    \I__879\ : InMux
    port map (
            O => \N__5005\,
            I => \N__4911\
        );

    \I__878\ : InMux
    port map (
            O => \N__5004\,
            I => \N__4900\
        );

    \I__877\ : InMux
    port map (
            O => \N__5003\,
            I => \N__4900\
        );

    \I__876\ : InMux
    port map (
            O => \N__5002\,
            I => \N__4900\
        );

    \I__875\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4900\
        );

    \I__874\ : InMux
    port map (
            O => \N__5000\,
            I => \N__4900\
        );

    \I__873\ : InMux
    port map (
            O => \N__4999\,
            I => \N__4885\
        );

    \I__872\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4885\
        );

    \I__871\ : InMux
    port map (
            O => \N__4997\,
            I => \N__4885\
        );

    \I__870\ : InMux
    port map (
            O => \N__4996\,
            I => \N__4885\
        );

    \I__869\ : InMux
    port map (
            O => \N__4995\,
            I => \N__4885\
        );

    \I__868\ : InMux
    port map (
            O => \N__4994\,
            I => \N__4885\
        );

    \I__867\ : InMux
    port map (
            O => \N__4993\,
            I => \N__4885\
        );

    \I__866\ : InMux
    port map (
            O => \N__4992\,
            I => \N__4868\
        );

    \I__865\ : InMux
    port map (
            O => \N__4991\,
            I => \N__4868\
        );

    \I__864\ : InMux
    port map (
            O => \N__4990\,
            I => \N__4868\
        );

    \I__863\ : InMux
    port map (
            O => \N__4989\,
            I => \N__4868\
        );

    \I__862\ : InMux
    port map (
            O => \N__4988\,
            I => \N__4868\
        );

    \I__861\ : InMux
    port map (
            O => \N__4987\,
            I => \N__4868\
        );

    \I__860\ : InMux
    port map (
            O => \N__4986\,
            I => \N__4868\
        );

    \I__859\ : InMux
    port map (
            O => \N__4985\,
            I => \N__4868\
        );

    \I__858\ : InMux
    port map (
            O => \N__4984\,
            I => \N__4847\
        );

    \I__857\ : InMux
    port map (
            O => \N__4983\,
            I => \N__4847\
        );

    \I__856\ : Span4Mux_s2_h
    port map (
            O => \N__4980\,
            I => \N__4842\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4973\,
            I => \N__4842\
        );

    \I__854\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4839\
        );

    \I__853\ : InMux
    port map (
            O => \N__4971\,
            I => \N__4828\
        );

    \I__852\ : InMux
    port map (
            O => \N__4970\,
            I => \N__4828\
        );

    \I__851\ : InMux
    port map (
            O => \N__4969\,
            I => \N__4828\
        );

    \I__850\ : InMux
    port map (
            O => \N__4968\,
            I => \N__4828\
        );

    \I__849\ : InMux
    port map (
            O => \N__4967\,
            I => \N__4828\
        );

    \I__848\ : InMux
    port map (
            O => \N__4966\,
            I => \N__4823\
        );

    \I__847\ : InMux
    port map (
            O => \N__4965\,
            I => \N__4823\
        );

    \I__846\ : InMux
    port map (
            O => \N__4964\,
            I => \N__4814\
        );

    \I__845\ : InMux
    port map (
            O => \N__4963\,
            I => \N__4814\
        );

    \I__844\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4814\
        );

    \I__843\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4814\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__4960\,
            I => \N__4811\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__4957\,
            I => \N__4803\
        );

    \I__840\ : InMux
    port map (
            O => \N__4956\,
            I => \N__4788\
        );

    \I__839\ : InMux
    port map (
            O => \N__4955\,
            I => \N__4788\
        );

    \I__838\ : InMux
    port map (
            O => \N__4954\,
            I => \N__4788\
        );

    \I__837\ : InMux
    port map (
            O => \N__4953\,
            I => \N__4788\
        );

    \I__836\ : InMux
    port map (
            O => \N__4952\,
            I => \N__4788\
        );

    \I__835\ : InMux
    port map (
            O => \N__4951\,
            I => \N__4788\
        );

    \I__834\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4788\
        );

    \I__833\ : InMux
    port map (
            O => \N__4949\,
            I => \N__4771\
        );

    \I__832\ : InMux
    port map (
            O => \N__4948\,
            I => \N__4771\
        );

    \I__831\ : InMux
    port map (
            O => \N__4947\,
            I => \N__4771\
        );

    \I__830\ : InMux
    port map (
            O => \N__4946\,
            I => \N__4771\
        );

    \I__829\ : InMux
    port map (
            O => \N__4945\,
            I => \N__4771\
        );

    \I__828\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4771\
        );

    \I__827\ : InMux
    port map (
            O => \N__4943\,
            I => \N__4771\
        );

    \I__826\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4771\
        );

    \I__825\ : Span4Mux_v
    port map (
            O => \N__4939\,
            I => \N__4756\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4932\,
            I => \N__4756\
        );

    \I__823\ : Span4Mux_h
    port map (
            O => \N__4927\,
            I => \N__4756\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4922\,
            I => \N__4756\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4911\,
            I => \N__4756\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__4900\,
            I => \N__4756\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__4885\,
            I => \N__4756\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__4868\,
            I => \N__4753\
        );

    \I__817\ : InMux
    port map (
            O => \N__4867\,
            I => \N__4738\
        );

    \I__816\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4738\
        );

    \I__815\ : InMux
    port map (
            O => \N__4865\,
            I => \N__4738\
        );

    \I__814\ : InMux
    port map (
            O => \N__4864\,
            I => \N__4738\
        );

    \I__813\ : InMux
    port map (
            O => \N__4863\,
            I => \N__4738\
        );

    \I__812\ : InMux
    port map (
            O => \N__4862\,
            I => \N__4738\
        );

    \I__811\ : InMux
    port map (
            O => \N__4861\,
            I => \N__4738\
        );

    \I__810\ : InMux
    port map (
            O => \N__4860\,
            I => \N__4721\
        );

    \I__809\ : InMux
    port map (
            O => \N__4859\,
            I => \N__4721\
        );

    \I__808\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4721\
        );

    \I__807\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4721\
        );

    \I__806\ : InMux
    port map (
            O => \N__4856\,
            I => \N__4721\
        );

    \I__805\ : InMux
    port map (
            O => \N__4855\,
            I => \N__4721\
        );

    \I__804\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4721\
        );

    \I__803\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4721\
        );

    \I__802\ : InMux
    port map (
            O => \N__4852\,
            I => \N__4718\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__4847\,
            I => \N__4707\
        );

    \I__800\ : Span4Mux_h
    port map (
            O => \N__4842\,
            I => \N__4707\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4839\,
            I => \N__4707\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4828\,
            I => \N__4707\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4823\,
            I => \N__4707\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__4814\,
            I => \N__4704\
        );

    \I__795\ : InMux
    port map (
            O => \N__4811\,
            I => \N__4701\
        );

    \I__794\ : CascadeMux
    port map (
            O => \N__4810\,
            I => \N__4698\
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__4809\,
            I => \N__4695\
        );

    \I__792\ : CascadeMux
    port map (
            O => \N__4808\,
            I => \N__4691\
        );

    \I__791\ : InMux
    port map (
            O => \N__4807\,
            I => \N__4684\
        );

    \I__790\ : InMux
    port map (
            O => \N__4806\,
            I => \N__4681\
        );

    \I__789\ : Span12Mux_s4_h
    port map (
            O => \N__4803\,
            I => \N__4674\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__4788\,
            I => \N__4674\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__4771\,
            I => \N__4674\
        );

    \I__786\ : Span4Mux_v
    port map (
            O => \N__4756\,
            I => \N__4665\
        );

    \I__785\ : Span4Mux_h
    port map (
            O => \N__4753\,
            I => \N__4665\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__4738\,
            I => \N__4665\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__4721\,
            I => \N__4665\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__4718\,
            I => \N__4656\
        );

    \I__781\ : Span4Mux_v
    port map (
            O => \N__4707\,
            I => \N__4656\
        );

    \I__780\ : Span4Mux_s2_h
    port map (
            O => \N__4704\,
            I => \N__4656\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__4701\,
            I => \N__4656\
        );

    \I__778\ : InMux
    port map (
            O => \N__4698\,
            I => \N__4651\
        );

    \I__777\ : InMux
    port map (
            O => \N__4695\,
            I => \N__4651\
        );

    \I__776\ : InMux
    port map (
            O => \N__4694\,
            I => \N__4648\
        );

    \I__775\ : InMux
    port map (
            O => \N__4691\,
            I => \N__4643\
        );

    \I__774\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4643\
        );

    \I__773\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4636\
        );

    \I__772\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4636\
        );

    \I__771\ : InMux
    port map (
            O => \N__4687\,
            I => \N__4636\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4684\,
            I => fsm_ctrl_inst1_current_state_1
        );

    \I__769\ : LocalMux
    port map (
            O => \N__4681\,
            I => fsm_ctrl_inst1_current_state_1
        );

    \I__768\ : Odrv12
    port map (
            O => \N__4674\,
            I => fsm_ctrl_inst1_current_state_1
        );

    \I__767\ : Odrv4
    port map (
            O => \N__4665\,
            I => fsm_ctrl_inst1_current_state_1
        );

    \I__766\ : Odrv4
    port map (
            O => \N__4656\,
            I => fsm_ctrl_inst1_current_state_1
        );

    \I__765\ : LocalMux
    port map (
            O => \N__4651\,
            I => fsm_ctrl_inst1_current_state_1
        );

    \I__764\ : LocalMux
    port map (
            O => \N__4648\,
            I => fsm_ctrl_inst1_current_state_1
        );

    \I__763\ : LocalMux
    port map (
            O => \N__4643\,
            I => fsm_ctrl_inst1_current_state_1
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4636\,
            I => fsm_ctrl_inst1_current_state_1
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__4617\,
            I => \config_register_latched_dec_inst1.STATSR_cnv_x1Z0Z_0_cascade_\
        );

    \I__760\ : InMux
    port map (
            O => \N__4614\,
            I => \N__4611\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__4611\,
            I => \config_register_latched_dec_inst1.STATSR_cnv_x0Z0Z_0\
        );

    \I__758\ : IoInMux
    port map (
            O => \N__4608\,
            I => \N__4605\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__4605\,
            I => \N__4602\
        );

    \I__756\ : Span12Mux_s11_v
    port map (
            O => \N__4602\,
            I => \N__4599\
        );

    \I__755\ : Odrv12
    port map (
            O => \N__4599\,
            I => \STATSR_cnv_ns_0\
        );

    \I__754\ : InMux
    port map (
            O => \N__4596\,
            I => \N__4585\
        );

    \I__753\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4570\
        );

    \I__752\ : InMux
    port map (
            O => \N__4594\,
            I => \N__4570\
        );

    \I__751\ : InMux
    port map (
            O => \N__4593\,
            I => \N__4570\
        );

    \I__750\ : InMux
    port map (
            O => \N__4592\,
            I => \N__4570\
        );

    \I__749\ : InMux
    port map (
            O => \N__4591\,
            I => \N__4570\
        );

    \I__748\ : InMux
    port map (
            O => \N__4590\,
            I => \N__4570\
        );

    \I__747\ : InMux
    port map (
            O => \N__4589\,
            I => \N__4560\
        );

    \I__746\ : InMux
    port map (
            O => \N__4588\,
            I => \N__4560\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__4585\,
            I => \N__4557\
        );

    \I__744\ : InMux
    port map (
            O => \N__4584\,
            I => \N__4536\
        );

    \I__743\ : InMux
    port map (
            O => \N__4583\,
            I => \N__4536\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4570\,
            I => \N__4533\
        );

    \I__741\ : InMux
    port map (
            O => \N__4569\,
            I => \N__4522\
        );

    \I__740\ : InMux
    port map (
            O => \N__4568\,
            I => \N__4522\
        );

    \I__739\ : InMux
    port map (
            O => \N__4567\,
            I => \N__4522\
        );

    \I__738\ : InMux
    port map (
            O => \N__4566\,
            I => \N__4522\
        );

    \I__737\ : InMux
    port map (
            O => \N__4565\,
            I => \N__4522\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__4560\,
            I => \N__4517\
        );

    \I__735\ : Span4Mux_s2_h
    port map (
            O => \N__4557\,
            I => \N__4517\
        );

    \I__734\ : InMux
    port map (
            O => \N__4556\,
            I => \N__4510\
        );

    \I__733\ : InMux
    port map (
            O => \N__4555\,
            I => \N__4510\
        );

    \I__732\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4510\
        );

    \I__731\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4504\
        );

    \I__730\ : InMux
    port map (
            O => \N__4552\,
            I => \N__4487\
        );

    \I__729\ : InMux
    port map (
            O => \N__4551\,
            I => \N__4487\
        );

    \I__728\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4487\
        );

    \I__727\ : InMux
    port map (
            O => \N__4549\,
            I => \N__4487\
        );

    \I__726\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4487\
        );

    \I__725\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4487\
        );

    \I__724\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4487\
        );

    \I__723\ : InMux
    port map (
            O => \N__4545\,
            I => \N__4487\
        );

    \I__722\ : InMux
    port map (
            O => \N__4544\,
            I => \N__4482\
        );

    \I__721\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4482\
        );

    \I__720\ : InMux
    port map (
            O => \N__4542\,
            I => \N__4477\
        );

    \I__719\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4477\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__4536\,
            I => \N__4466\
        );

    \I__717\ : Span4Mux_v
    port map (
            O => \N__4533\,
            I => \N__4466\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__4522\,
            I => \N__4466\
        );

    \I__715\ : Span4Mux_v
    port map (
            O => \N__4517\,
            I => \N__4466\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__4510\,
            I => \N__4466\
        );

    \I__713\ : InMux
    port map (
            O => \N__4509\,
            I => \N__4459\
        );

    \I__712\ : InMux
    port map (
            O => \N__4508\,
            I => \N__4459\
        );

    \I__711\ : InMux
    port map (
            O => \N__4507\,
            I => \N__4459\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4504\,
            I => fsm_ctrl_inst1_current_state_0
        );

    \I__709\ : LocalMux
    port map (
            O => \N__4487\,
            I => fsm_ctrl_inst1_current_state_0
        );

    \I__708\ : LocalMux
    port map (
            O => \N__4482\,
            I => fsm_ctrl_inst1_current_state_0
        );

    \I__707\ : LocalMux
    port map (
            O => \N__4477\,
            I => fsm_ctrl_inst1_current_state_0
        );

    \I__706\ : Odrv4
    port map (
            O => \N__4466\,
            I => fsm_ctrl_inst1_current_state_0
        );

    \I__705\ : LocalMux
    port map (
            O => \N__4459\,
            I => fsm_ctrl_inst1_current_state_0
        );

    \I__704\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4443\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__4443\,
            I => \N__4436\
        );

    \I__702\ : InMux
    port map (
            O => \N__4442\,
            I => \N__4429\
        );

    \I__701\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4429\
        );

    \I__700\ : InMux
    port map (
            O => \N__4440\,
            I => \N__4429\
        );

    \I__699\ : InMux
    port map (
            O => \N__4439\,
            I => \N__4426\
        );

    \I__698\ : Odrv4
    port map (
            O => \N__4436\,
            I => \SEL_REG\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__4429\,
            I => \SEL_REG\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__4426\,
            I => \SEL_REG\
        );

    \I__695\ : InMux
    port map (
            O => \N__4419\,
            I => \N__4415\
        );

    \I__694\ : InMux
    port map (
            O => \N__4418\,
            I => \N__4412\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__4415\,
            I => \N__4409\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__4412\,
            I => \MOSI\
        );

    \I__691\ : Odrv4
    port map (
            O => \N__4409\,
            I => \MOSI\
        );

    \I__690\ : InMux
    port map (
            O => \N__4404\,
            I => \N__4401\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__4401\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_0\
        );

    \I__688\ : InMux
    port map (
            O => \N__4398\,
            I => \N__4395\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__4395\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_1\
        );

    \I__686\ : InMux
    port map (
            O => \N__4392\,
            I => \N__4389\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4389\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_2\
        );

    \I__684\ : InMux
    port map (
            O => \N__4386\,
            I => \N__4383\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__4383\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_3\
        );

    \I__682\ : InMux
    port map (
            O => \N__4380\,
            I => \N__4377\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4377\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_1\
        );

    \I__680\ : InMux
    port map (
            O => \N__4374\,
            I => \N__4371\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__4371\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_14\
        );

    \I__678\ : InMux
    port map (
            O => \N__4368\,
            I => \N__4365\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4365\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_15\
        );

    \I__676\ : InMux
    port map (
            O => \N__4362\,
            I => \N__4359\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__4359\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_12\
        );

    \I__674\ : InMux
    port map (
            O => \N__4356\,
            I => \N__4353\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__4353\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_13\
        );

    \I__672\ : InMux
    port map (
            O => \N__4350\,
            I => \N__4347\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4347\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_10\
        );

    \I__670\ : InMux
    port map (
            O => \N__4344\,
            I => \N__4341\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__4341\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_11\
        );

    \I__668\ : CascadeMux
    port map (
            O => \N__4338\,
            I => \config_register_latched_dec_inst1.DYNSR_cnv_x0Z0Z_0_cascade_\
        );

    \I__667\ : InMux
    port map (
            O => \N__4335\,
            I => \N__4332\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__4332\,
            I => \config_register_latched_dec_inst1.DYNSR_cnv_x1Z0Z_0\
        );

    \I__665\ : InMux
    port map (
            O => \N__4329\,
            I => \N__4317\
        );

    \I__664\ : InMux
    port map (
            O => \N__4328\,
            I => \N__4317\
        );

    \I__663\ : InMux
    port map (
            O => \N__4327\,
            I => \N__4317\
        );

    \I__662\ : InMux
    port map (
            O => \N__4326\,
            I => \N__4317\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4317\,
            I => \fsm_ctrl_inst1.counter_dinZ0Z_2\
        );

    \I__660\ : CascadeMux
    port map (
            O => \N__4314\,
            I => \N__4309\
        );

    \I__659\ : CascadeMux
    port map (
            O => \N__4313\,
            I => \N__4306\
        );

    \I__658\ : CascadeMux
    port map (
            O => \N__4312\,
            I => \N__4303\
        );

    \I__657\ : InMux
    port map (
            O => \N__4309\,
            I => \N__4296\
        );

    \I__656\ : InMux
    port map (
            O => \N__4306\,
            I => \N__4296\
        );

    \I__655\ : InMux
    port map (
            O => \N__4303\,
            I => \N__4296\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4296\,
            I => \fsm_ctrl_inst1.counter_dinZ0Z_3\
        );

    \I__653\ : CascadeMux
    port map (
            O => \N__4293\,
            I => \N__4289\
        );

    \I__652\ : InMux
    port map (
            O => \N__4292\,
            I => \N__4275\
        );

    \I__651\ : InMux
    port map (
            O => \N__4289\,
            I => \N__4275\
        );

    \I__650\ : InMux
    port map (
            O => \N__4288\,
            I => \N__4275\
        );

    \I__649\ : InMux
    port map (
            O => \N__4287\,
            I => \N__4275\
        );

    \I__648\ : InMux
    port map (
            O => \N__4286\,
            I => \N__4275\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__4275\,
            I => \fsm_ctrl_inst1.counter_dinZ0Z_1\
        );

    \I__646\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4264\
        );

    \I__645\ : InMux
    port map (
            O => \N__4271\,
            I => \N__4255\
        );

    \I__644\ : InMux
    port map (
            O => \N__4270\,
            I => \N__4255\
        );

    \I__643\ : InMux
    port map (
            O => \N__4269\,
            I => \N__4255\
        );

    \I__642\ : InMux
    port map (
            O => \N__4268\,
            I => \N__4255\
        );

    \I__641\ : InMux
    port map (
            O => \N__4267\,
            I => \N__4252\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__4264\,
            I => \N__4247\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4255\,
            I => \N__4247\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__4252\,
            I => \fsm_ctrl_inst1.counter_dinZ0Z_0\
        );

    \I__637\ : Odrv4
    port map (
            O => \N__4247\,
            I => \fsm_ctrl_inst1.counter_dinZ0Z_0\
        );

    \I__636\ : CascadeMux
    port map (
            O => \N__4242\,
            I => \fsm_ctrl_inst1.o2_cascade_\
        );

    \I__635\ : InMux
    port map (
            O => \N__4239\,
            I => \N__4236\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__4236\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_0\
        );

    \I__633\ : InMux
    port map (
            O => \N__4233\,
            I => \N__4230\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__4230\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_19\
        );

    \I__631\ : InMux
    port map (
            O => \N__4227\,
            I => \N__4224\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4224\,
            I => \N__4221\
        );

    \I__629\ : Odrv4
    port map (
            O => \N__4221\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_20\
        );

    \I__628\ : CEMux
    port map (
            O => \N__4218\,
            I => \N__4155\
        );

    \I__627\ : CEMux
    port map (
            O => \N__4217\,
            I => \N__4155\
        );

    \I__626\ : CEMux
    port map (
            O => \N__4216\,
            I => \N__4155\
        );

    \I__625\ : CEMux
    port map (
            O => \N__4215\,
            I => \N__4155\
        );

    \I__624\ : CEMux
    port map (
            O => \N__4214\,
            I => \N__4155\
        );

    \I__623\ : CEMux
    port map (
            O => \N__4213\,
            I => \N__4155\
        );

    \I__622\ : CEMux
    port map (
            O => \N__4212\,
            I => \N__4155\
        );

    \I__621\ : CEMux
    port map (
            O => \N__4211\,
            I => \N__4155\
        );

    \I__620\ : CEMux
    port map (
            O => \N__4210\,
            I => \N__4155\
        );

    \I__619\ : CEMux
    port map (
            O => \N__4209\,
            I => \N__4155\
        );

    \I__618\ : CEMux
    port map (
            O => \N__4208\,
            I => \N__4155\
        );

    \I__617\ : CEMux
    port map (
            O => \N__4207\,
            I => \N__4155\
        );

    \I__616\ : CEMux
    port map (
            O => \N__4206\,
            I => \N__4155\
        );

    \I__615\ : CEMux
    port map (
            O => \N__4205\,
            I => \N__4155\
        );

    \I__614\ : CEMux
    port map (
            O => \N__4204\,
            I => \N__4155\
        );

    \I__613\ : CEMux
    port map (
            O => \N__4203\,
            I => \N__4155\
        );

    \I__612\ : CEMux
    port map (
            O => \N__4202\,
            I => \N__4155\
        );

    \I__611\ : CEMux
    port map (
            O => \N__4201\,
            I => \N__4155\
        );

    \I__610\ : CEMux
    port map (
            O => \N__4200\,
            I => \N__4155\
        );

    \I__609\ : CEMux
    port map (
            O => \N__4199\,
            I => \N__4155\
        );

    \I__608\ : CEMux
    port map (
            O => \N__4198\,
            I => \N__4155\
        );

    \I__607\ : GlobalMux
    port map (
            O => \N__4155\,
            I => \N__4152\
        );

    \I__606\ : gio2CtrlBuf
    port map (
            O => \N__4152\,
            I => \fsm_ctrl_inst1.current_state_i_g_0\
        );

    \I__605\ : IoInMux
    port map (
            O => \N__4149\,
            I => \N__4146\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__4146\,
            I => \N__4143\
        );

    \I__603\ : IoSpan4Mux
    port map (
            O => \N__4143\,
            I => \N__4140\
        );

    \I__602\ : Span4Mux_s3_h
    port map (
            O => \N__4140\,
            I => \N__4137\
        );

    \I__601\ : Odrv4
    port map (
            O => \N__4137\,
            I => \SDO_signal_out_c\
        );

    \I__600\ : InMux
    port map (
            O => \N__4134\,
            I => \N__4131\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__4131\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_31\
        );

    \I__598\ : InMux
    port map (
            O => \N__4128\,
            I => \N__4125\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__4125\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_32\
        );

    \I__596\ : InMux
    port map (
            O => \N__4122\,
            I => \N__4109\
        );

    \I__595\ : InMux
    port map (
            O => \N__4121\,
            I => \N__4109\
        );

    \I__594\ : InMux
    port map (
            O => \N__4120\,
            I => \N__4109\
        );

    \I__593\ : InMux
    port map (
            O => \N__4119\,
            I => \N__4106\
        );

    \I__592\ : InMux
    port map (
            O => \N__4118\,
            I => \N__4103\
        );

    \I__591\ : InMux
    port map (
            O => \N__4117\,
            I => \N__4100\
        );

    \I__590\ : InMux
    port map (
            O => \N__4116\,
            I => \N__4097\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__4109\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_1\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__4106\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_1\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4103\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_1\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4100\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_1\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__4097\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_1\
        );

    \I__584\ : CascadeMux
    port map (
            O => \N__4086\,
            I => \N__4081\
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__4085\,
            I => \N__4078\
        );

    \I__582\ : InMux
    port map (
            O => \N__4084\,
            I => \N__4071\
        );

    \I__581\ : InMux
    port map (
            O => \N__4081\,
            I => \N__4064\
        );

    \I__580\ : InMux
    port map (
            O => \N__4078\,
            I => \N__4064\
        );

    \I__579\ : InMux
    port map (
            O => \N__4077\,
            I => \N__4064\
        );

    \I__578\ : InMux
    port map (
            O => \N__4076\,
            I => \N__4061\
        );

    \I__577\ : InMux
    port map (
            O => \N__4075\,
            I => \N__4058\
        );

    \I__576\ : InMux
    port map (
            O => \N__4074\,
            I => \N__4055\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__4071\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_3\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__4064\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_3\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4061\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_3\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4058\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_3\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4055\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_3\
        );

    \I__570\ : InMux
    port map (
            O => \N__4044\,
            I => \N__4039\
        );

    \I__569\ : InMux
    port map (
            O => \N__4043\,
            I => \N__4036\
        );

    \I__568\ : InMux
    port map (
            O => \N__4042\,
            I => \N__4033\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4039\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_0\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4036\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_0\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__4033\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_0\
        );

    \I__564\ : InMux
    port map (
            O => \N__4026\,
            I => \N__4023\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4023\,
            I => \fsm_ctrl_inst1.current_state_RNO_2Z0Z_0\
        );

    \I__562\ : InMux
    port map (
            O => \N__4020\,
            I => \N__4017\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__4017\,
            I => \fsm_ctrl_inst1.g0_0_3_0\
        );

    \I__560\ : CascadeMux
    port map (
            O => \N__4014\,
            I => \N__4007\
        );

    \I__559\ : CascadeMux
    port map (
            O => \N__4013\,
            I => \N__4002\
        );

    \I__558\ : InMux
    port map (
            O => \N__4012\,
            I => \N__3999\
        );

    \I__557\ : InMux
    port map (
            O => \N__4011\,
            I => \N__3996\
        );

    \I__556\ : InMux
    port map (
            O => \N__4010\,
            I => \N__3993\
        );

    \I__555\ : InMux
    port map (
            O => \N__4007\,
            I => \N__3990\
        );

    \I__554\ : InMux
    port map (
            O => \N__4006\,
            I => \N__3983\
        );

    \I__553\ : InMux
    port map (
            O => \N__4005\,
            I => \N__3983\
        );

    \I__552\ : InMux
    port map (
            O => \N__4002\,
            I => \N__3983\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3999\,
            I => \fsm_ctrl_inst1.counter_idleZ1Z_4\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__3996\,
            I => \fsm_ctrl_inst1.counter_idleZ1Z_4\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3993\,
            I => \fsm_ctrl_inst1.counter_idleZ1Z_4\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3990\,
            I => \fsm_ctrl_inst1.counter_idleZ1Z_4\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3983\,
            I => \fsm_ctrl_inst1.counter_idleZ1Z_4\
        );

    \I__546\ : InMux
    port map (
            O => \N__3972\,
            I => \N__3963\
        );

    \I__545\ : InMux
    port map (
            O => \N__3971\,
            I => \N__3958\
        );

    \I__544\ : InMux
    port map (
            O => \N__3970\,
            I => \N__3958\
        );

    \I__543\ : InMux
    port map (
            O => \N__3969\,
            I => \N__3955\
        );

    \I__542\ : InMux
    port map (
            O => \N__3968\,
            I => \N__3950\
        );

    \I__541\ : InMux
    port map (
            O => \N__3967\,
            I => \N__3950\
        );

    \I__540\ : InMux
    port map (
            O => \N__3966\,
            I => \N__3947\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3963\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_2\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3958\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_2\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3955\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_2\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3950\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_2\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3947\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_2\
        );

    \I__534\ : InMux
    port map (
            O => \N__3936\,
            I => \N__3933\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3933\,
            I => \fsm_ctrl_inst1.g0_0_3\
        );

    \I__532\ : CascadeMux
    port map (
            O => \N__3930\,
            I => \fsm_ctrl_inst1.counter_din_RNO_0Z0Z_3_cascade_\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__3927\,
            I => \fsm_ctrl_inst1.current_state_RNO_3Z0Z_0_cascade_\
        );

    \I__530\ : InMux
    port map (
            O => \N__3924\,
            I => \N__3921\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__3921\,
            I => \fsm_ctrl_inst1.current_state_RNO_1Z0Z_0\
        );

    \I__528\ : InMux
    port map (
            O => \N__3918\,
            I => \N__3915\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3915\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_23\
        );

    \I__526\ : InMux
    port map (
            O => \N__3912\,
            I => \N__3909\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3909\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_24\
        );

    \I__524\ : InMux
    port map (
            O => \N__3906\,
            I => \N__3903\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__3903\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_45\
        );

    \I__522\ : InMux
    port map (
            O => \N__3900\,
            I => \N__3897\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3897\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_46\
        );

    \I__520\ : InMux
    port map (
            O => \N__3894\,
            I => \N__3891\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3891\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_27\
        );

    \I__518\ : InMux
    port map (
            O => \N__3888\,
            I => \N__3885\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3885\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_28\
        );

    \I__516\ : InMux
    port map (
            O => \N__3882\,
            I => \N__3879\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3879\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_33\
        );

    \I__514\ : InMux
    port map (
            O => \N__3876\,
            I => \N__3873\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3873\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_29\
        );

    \I__512\ : InMux
    port map (
            O => \N__3870\,
            I => \N__3867\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3867\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_34\
        );

    \I__510\ : InMux
    port map (
            O => \N__3864\,
            I => \N__3861\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3861\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_30\
        );

    \I__508\ : InMux
    port map (
            O => \N__3858\,
            I => \N__3855\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3855\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_35\
        );

    \I__506\ : InMux
    port map (
            O => \N__3852\,
            I => \N__3849\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3849\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_36\
        );

    \I__504\ : InMux
    port map (
            O => \N__3846\,
            I => \N__3843\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3843\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_26\
        );

    \I__502\ : InMux
    port map (
            O => \N__3840\,
            I => \N__3837\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__3837\,
            I => \N__3834\
        );

    \I__500\ : Odrv4
    port map (
            O => \N__3834\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_12\
        );

    \I__499\ : InMux
    port map (
            O => \N__3831\,
            I => \N__3828\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3828\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_13\
        );

    \I__497\ : InMux
    port map (
            O => \N__3825\,
            I => \N__3822\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__3822\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_49\
        );

    \I__495\ : InMux
    port map (
            O => \N__3819\,
            I => \N__3816\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3816\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_50\
        );

    \I__493\ : InMux
    port map (
            O => \N__3813\,
            I => \N__3810\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3810\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_47\
        );

    \I__491\ : InMux
    port map (
            O => \N__3807\,
            I => \N__3804\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3804\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_25\
        );

    \I__489\ : InMux
    port map (
            O => \N__3801\,
            I => \N__3798\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__3798\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_44\
        );

    \I__487\ : InMux
    port map (
            O => \N__3795\,
            I => \N__3792\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3792\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_51\
        );

    \I__485\ : InMux
    port map (
            O => \N__3789\,
            I => \N__3786\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3786\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_52\
        );

    \I__483\ : InMux
    port map (
            O => \N__3783\,
            I => \N__3780\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3780\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_17\
        );

    \I__481\ : InMux
    port map (
            O => \N__3777\,
            I => \N__3774\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3774\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_16\
        );

    \I__479\ : InMux
    port map (
            O => \N__3771\,
            I => \N__3768\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__3768\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_14\
        );

    \I__477\ : InMux
    port map (
            O => \N__3765\,
            I => \N__3762\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3762\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_15\
        );

    \I__475\ : InMux
    port map (
            O => \N__3759\,
            I => \N__3756\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__3756\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_62\
        );

    \I__473\ : InMux
    port map (
            O => \N__3753\,
            I => \N__3750\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__3750\,
            I => \N__3747\
        );

    \I__471\ : Odrv12
    port map (
            O => \N__3747\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_63\
        );

    \I__470\ : InMux
    port map (
            O => \N__3744\,
            I => \N__3741\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3741\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_21\
        );

    \I__468\ : InMux
    port map (
            O => \N__3738\,
            I => \N__3735\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__3735\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_22\
        );

    \I__466\ : InMux
    port map (
            O => \N__3732\,
            I => \N__3729\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3729\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_48\
        );

    \I__464\ : InMux
    port map (
            O => \N__3726\,
            I => \N__3723\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__3723\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_65\
        );

    \I__462\ : InMux
    port map (
            O => \N__3720\,
            I => \N__3717\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__3717\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_66\
        );

    \I__460\ : InMux
    port map (
            O => \N__3714\,
            I => \N__3711\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3711\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_68\
        );

    \I__458\ : InMux
    port map (
            O => \N__3708\,
            I => \N__3705\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3705\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_69\
        );

    \I__456\ : InMux
    port map (
            O => \N__3702\,
            I => \N__3699\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__3699\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_70\
        );

    \I__454\ : InMux
    port map (
            O => \N__3696\,
            I => \N__3693\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3693\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_73\
        );

    \I__452\ : InMux
    port map (
            O => \N__3690\,
            I => \N__3687\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__3687\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_74\
        );

    \I__450\ : InMux
    port map (
            O => \N__3684\,
            I => \N__3681\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__3681\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_71\
        );

    \I__448\ : InMux
    port map (
            O => \N__3678\,
            I => \N__3675\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__3675\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_72\
        );

    \I__446\ : InMux
    port map (
            O => \N__3672\,
            I => \N__3669\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__3669\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_18\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__3666\,
            I => \fsm_ctrl_inst1.counter_idle_RNO_1Z0Z_0_cascade_\
        );

    \I__443\ : CascadeMux
    port map (
            O => \N__3663\,
            I => \fsm_ctrl_inst1.counter_idlee_0_cascade_\
        );

    \I__442\ : InMux
    port map (
            O => \N__3660\,
            I => \N__3657\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3657\,
            I => \fsm_ctrl_inst1.counter_idle_s_1\
        );

    \I__440\ : InMux
    port map (
            O => \N__3654\,
            I => \N__3651\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__3651\,
            I => \fsm_ctrl_inst1.g0_0_3_2\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__3648\,
            I => \N__3645\
        );

    \I__437\ : InMux
    port map (
            O => \N__3645\,
            I => \N__3642\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3642\,
            I => \fsm_ctrl_inst1.g0_0_2_2\
        );

    \I__435\ : InMux
    port map (
            O => \N__3639\,
            I => \N__3631\
        );

    \I__434\ : InMux
    port map (
            O => \N__3638\,
            I => \N__3631\
        );

    \I__433\ : InMux
    port map (
            O => \N__3637\,
            I => \N__3626\
        );

    \I__432\ : InMux
    port map (
            O => \N__3636\,
            I => \N__3626\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__3631\,
            I => \fsm_ctrl_inst1.current_state_20_d_i\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__3626\,
            I => \fsm_ctrl_inst1.current_state_20_d_i\
        );

    \I__429\ : InMux
    port map (
            O => \N__3621\,
            I => \N__3618\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3618\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_15\
        );

    \I__427\ : CascadeMux
    port map (
            O => \N__3615\,
            I => \N__3612\
        );

    \I__426\ : InMux
    port map (
            O => \N__3612\,
            I => \N__3609\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__3609\,
            I => \N__3606\
        );

    \I__424\ : Span4Mux_v
    port map (
            O => \N__3606\,
            I => \N__3603\
        );

    \I__423\ : Odrv4
    port map (
            O => \N__3603\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_87\
        );

    \I__422\ : InMux
    port map (
            O => \N__3600\,
            I => \N__3597\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3597\,
            I => \N__3594\
        );

    \I__420\ : Odrv4
    port map (
            O => \N__3594\,
            I => \CONSTANT_ONE_NET\
        );

    \I__419\ : InMux
    port map (
            O => \N__3591\,
            I => \N__3588\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__3588\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_67\
        );

    \I__417\ : InMux
    port map (
            O => \N__3585\,
            I => \N__3582\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__3582\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_64\
        );

    \I__415\ : CascadeMux
    port map (
            O => \N__3579\,
            I => \fsm_ctrl_inst1.g0_0_2_0_cascade_\
        );

    \I__414\ : InMux
    port map (
            O => \N__3576\,
            I => \N__3573\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__3573\,
            I => \fsm_ctrl_inst1.counter_idle_s_3\
        );

    \I__412\ : CascadeMux
    port map (
            O => \N__3570\,
            I => \fsm_ctrl_inst1.g0_0_2_cascade_\
        );

    \I__411\ : InMux
    port map (
            O => \N__3567\,
            I => \N__3564\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__3564\,
            I => \fsm_ctrl_inst1.counter_idle_s_4\
        );

    \I__409\ : InMux
    port map (
            O => \N__3561\,
            I => \N__3558\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__3558\,
            I => \fsm_ctrl_inst1.g0_0_3_1\
        );

    \I__407\ : InMux
    port map (
            O => \N__3555\,
            I => \N__3552\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__3552\,
            I => \fsm_ctrl_inst1.g0_0_2_1\
        );

    \I__405\ : CascadeMux
    port map (
            O => \N__3549\,
            I => \fsm_ctrl_inst1.current_state_20_d_i_cascade_\
        );

    \I__404\ : InMux
    port map (
            O => \N__3546\,
            I => \N__3543\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__3543\,
            I => \fsm_ctrl_inst1.counter_idle_s_2\
        );

    \I__402\ : CascadeMux
    port map (
            O => \N__3540\,
            I => \fsm_ctrl_inst1.N_93_0_cascade_\
        );

    \I__401\ : InMux
    port map (
            O => \N__3537\,
            I => \N__3534\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__3534\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_3\
        );

    \I__399\ : InMux
    port map (
            O => \N__3531\,
            I => \N__3528\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__3528\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_1\
        );

    \I__397\ : InMux
    port map (
            O => \N__3525\,
            I => \N__3522\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__3522\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_2\
        );

    \I__395\ : InMux
    port map (
            O => \N__3519\,
            I => \N__3516\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3516\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_38\
        );

    \I__393\ : InMux
    port map (
            O => \N__3513\,
            I => \N__3510\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__3510\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_39\
        );

    \I__391\ : InMux
    port map (
            O => \N__3507\,
            I => \N__3504\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3504\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_0\
        );

    \I__389\ : InMux
    port map (
            O => \N__3501\,
            I => \N__3498\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__3498\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_40\
        );

    \I__387\ : InMux
    port map (
            O => \N__3495\,
            I => \N__3492\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__3492\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_41\
        );

    \I__385\ : InMux
    port map (
            O => \N__3489\,
            I => \N__3486\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__3486\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_43\
        );

    \I__383\ : InMux
    port map (
            O => \N__3483\,
            I => \N__3480\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3480\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_80\
        );

    \I__381\ : InMux
    port map (
            O => \N__3477\,
            I => \N__3474\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__3474\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_4\
        );

    \I__379\ : InMux
    port map (
            O => \N__3471\,
            I => \N__3468\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__3468\,
            I => \N__3465\
        );

    \I__377\ : Odrv12
    port map (
            O => \N__3465\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_5\
        );

    \I__376\ : InMux
    port map (
            O => \N__3462\,
            I => \N__3459\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__3459\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_53\
        );

    \I__374\ : InMux
    port map (
            O => \N__3456\,
            I => \N__3453\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__3453\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_37\
        );

    \I__372\ : InMux
    port map (
            O => \N__3450\,
            I => \N__3447\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__3447\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_81\
        );

    \I__370\ : InMux
    port map (
            O => \N__3444\,
            I => \N__3441\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__3441\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_82\
        );

    \I__368\ : InMux
    port map (
            O => \N__3438\,
            I => \N__3435\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__3435\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_75\
        );

    \I__366\ : InMux
    port map (
            O => \N__3432\,
            I => \N__3429\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__3429\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_76\
        );

    \I__364\ : InMux
    port map (
            O => \N__3426\,
            I => \N__3423\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__3423\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_77\
        );

    \I__362\ : InMux
    port map (
            O => \N__3420\,
            I => \N__3417\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__3417\,
            I => \N__3414\
        );

    \I__360\ : Odrv4
    port map (
            O => \N__3414\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_11\
        );

    \I__359\ : InMux
    port map (
            O => \N__3411\,
            I => \N__3408\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3408\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_54\
        );

    \I__357\ : InMux
    port map (
            O => \N__3405\,
            I => \N__3402\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__3402\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_60\
        );

    \I__355\ : InMux
    port map (
            O => \N__3399\,
            I => \N__3396\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__3396\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_61\
        );

    \I__353\ : InMux
    port map (
            O => \N__3393\,
            I => \N__3390\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__3390\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_78\
        );

    \I__351\ : InMux
    port map (
            O => \N__3387\,
            I => \N__3384\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__3384\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_79\
        );

    \I__349\ : InMux
    port map (
            O => \N__3381\,
            I => \N__3378\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__3378\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_9\
        );

    \I__347\ : InMux
    port map (
            O => \N__3375\,
            I => \N__3372\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__3372\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_6\
        );

    \I__345\ : InMux
    port map (
            O => \N__3369\,
            I => \N__3366\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__3366\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_7\
        );

    \I__343\ : InMux
    port map (
            O => \N__3363\,
            I => \N__3360\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__3360\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_8\
        );

    \I__341\ : InMux
    port map (
            O => \N__3357\,
            I => \N__3354\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__3354\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_12\
        );

    \I__339\ : InMux
    port map (
            O => \N__3351\,
            I => \N__3348\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__3348\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_10\
        );

    \I__337\ : InMux
    port map (
            O => \N__3345\,
            I => \N__3342\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__3342\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_11\
        );

    \I__335\ : InMux
    port map (
            O => \N__3339\,
            I => \N__3336\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__3336\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_13\
        );

    \I__333\ : InMux
    port map (
            O => \N__3333\,
            I => \N__3330\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__3330\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_14\
        );

    \I__331\ : CEMux
    port map (
            O => \N__3327\,
            I => \N__3322\
        );

    \I__330\ : CEMux
    port map (
            O => \N__3326\,
            I => \N__3319\
        );

    \I__329\ : CEMux
    port map (
            O => \N__3325\,
            I => \N__3316\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__3322\,
            I => \N__3313\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__3319\,
            I => \N__3308\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__3316\,
            I => \N__3308\
        );

    \I__325\ : Odrv4
    port map (
            O => \N__3313\,
            I => \fsm_ctrl_inst1.current_state_i_1\
        );

    \I__324\ : Odrv4
    port map (
            O => \N__3308\,
            I => \fsm_ctrl_inst1.current_state_i_1\
        );

    \I__323\ : InMux
    port map (
            O => \N__3303\,
            I => \N__3300\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__3300\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_42\
        );

    \I__321\ : InMux
    port map (
            O => \N__3297\,
            I => \fsm_ctrl_inst1.counter_idle_cry_0\
        );

    \I__320\ : InMux
    port map (
            O => \N__3294\,
            I => \fsm_ctrl_inst1.counter_idle_cry_1\
        );

    \I__319\ : InMux
    port map (
            O => \N__3291\,
            I => \fsm_ctrl_inst1.counter_idle_cry_2\
        );

    \I__318\ : InMux
    port map (
            O => \N__3288\,
            I => \fsm_ctrl_inst1.counter_idle_cry_3\
        );

    \I__317\ : InMux
    port map (
            O => \N__3285\,
            I => \N__3282\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__3282\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_3\
        );

    \I__315\ : InMux
    port map (
            O => \N__3279\,
            I => \N__3276\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__3276\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_4\
        );

    \I__313\ : InMux
    port map (
            O => \N__3273\,
            I => \N__3270\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__3270\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_56\
        );

    \I__311\ : InMux
    port map (
            O => \N__3267\,
            I => \N__3264\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__3264\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_59\
        );

    \I__309\ : InMux
    port map (
            O => \N__3261\,
            I => \N__3258\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__3258\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_55\
        );

    \I__307\ : InMux
    port map (
            O => \N__3255\,
            I => \N__3252\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__3252\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_7\
        );

    \I__305\ : InMux
    port map (
            O => \N__3249\,
            I => \N__3246\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__3246\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_8\
        );

    \I__303\ : InMux
    port map (
            O => \N__3243\,
            I => \N__3240\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__3240\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_9\
        );

    \I__301\ : InMux
    port map (
            O => \N__3237\,
            I => \N__3234\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__3234\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_10\
        );

    \I__299\ : InMux
    port map (
            O => \N__3231\,
            I => \N__3228\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__3228\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_83\
        );

    \I__297\ : InMux
    port map (
            O => \N__3225\,
            I => \N__3222\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__3222\,
            I => \N__3219\
        );

    \I__295\ : Odrv4
    port map (
            O => \N__3219\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_84\
        );

    \I__294\ : InMux
    port map (
            O => \N__3216\,
            I => \N__3213\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__3213\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_85\
        );

    \I__292\ : InMux
    port map (
            O => \N__3210\,
            I => \N__3207\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__3207\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_86\
        );

    \I__290\ : InMux
    port map (
            O => \N__3204\,
            I => \N__3201\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__3201\,
            I => \N__3198\
        );

    \I__288\ : Odrv4
    port map (
            O => \N__3198\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_1\
        );

    \I__287\ : InMux
    port map (
            O => \N__3195\,
            I => \N__3192\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__3192\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_2\
        );

    \I__285\ : InMux
    port map (
            O => \N__3189\,
            I => \N__3186\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__3186\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_5\
        );

    \I__283\ : InMux
    port map (
            O => \N__3183\,
            I => \N__3180\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__3180\,
            I => \N__3177\
        );

    \I__281\ : Span4Mux_v
    port map (
            O => \N__3177\,
            I => \N__3174\
        );

    \I__280\ : Odrv4
    port map (
            O => \N__3174\,
            I => \RST_N_c\
        );

    \I__279\ : IoInMux
    port map (
            O => \N__3171\,
            I => \N__3168\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__3168\,
            I => \N__3165\
        );

    \I__277\ : Span12Mux_s0_h
    port map (
            O => \N__3165\,
            I => \N__3162\
        );

    \I__276\ : Odrv12
    port map (
            O => \N__3162\,
            I => \RST_N_c_i\
        );

    \I__275\ : IoInMux
    port map (
            O => \N__3159\,
            I => \N__3156\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__3156\,
            I => \fsm_ctrl_inst1.current_state_i_0\
        );

    \I__273\ : InMux
    port map (
            O => \N__3153\,
            I => \N__3150\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__3150\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_58\
        );

    \I__271\ : InMux
    port map (
            O => \N__3147\,
            I => \N__3144\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__3144\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_57\
        );

    \I__269\ : InMux
    port map (
            O => \N__3141\,
            I => \N__3138\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__3138\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_6\
        );

    \I__267\ : InMux
    port map (
            O => \N__3135\,
            I => \N__3132\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__3132\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_0\
        );

    \IN_MUX_bfv_3_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_20_0_\
        );

    \N_218_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4608\,
            GLOBALBUFFEROUTPUT => \N_218_g\
        );

    \fsm_ctrl_inst1.current_state_RNI1GR8_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3159\,
            GLOBALBUFFEROUTPUT => \fsm_ctrl_inst1.current_state_i_g_0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \RST_N_ibuf_RNIBJGC_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3171\,
            GLOBALBUFFEROUTPUT => \RST_N_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \RST_N_ibuf_RNIBJGC_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3183\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RST_N_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.current_state_RNI1GR8_0_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4596\,
            lcout => \fsm_ctrl_inst1.current_state_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_58_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3147\,
            in2 => \_gnd_net_\,
            in3 => \N__5036\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6121\,
            ce => \N__4200\,
            sr => \N__5801\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_59_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5055\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3153\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6119\,
            ce => \N__4198\,
            sr => \N__5802\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_57_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3273\,
            in2 => \_gnd_net_\,
            in3 => \N__5054\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6119\,
            ce => \N__4198\,
            sr => \N__5802\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_7_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3141\,
            in2 => \_gnd_net_\,
            in3 => \N__4984\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6122\,
            ce => \N__4201\,
            sr => \N__5804\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_6_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3471\,
            in2 => \_gnd_net_\,
            in3 => \N__4983\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6122\,
            ce => \N__4201\,
            sr => \N__5804\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_84_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3231\,
            in2 => \_gnd_net_\,
            in3 => \N__4972\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6124\,
            ce => \N__4203\,
            sr => \N__5807\
        );

    \fsm_ctrl_inst1.bit_sequence_din_1_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4588\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3135\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6127\,
            ce => \N__3325\,
            sr => \N__5811\
        );

    \fsm_ctrl_inst1.bit_sequence_din_0_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4589\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6127\,
            ce => \N__3325\,
            sr => \N__5811\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_85_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3225\,
            in2 => \_gnd_net_\,
            in3 => \N__4962\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6131\,
            ce => \N__4209\,
            sr => \N__5816\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_86_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4963\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3216\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6131\,
            ce => \N__4209\,
            sr => \N__5816\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_87_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3210\,
            in2 => \_gnd_net_\,
            in3 => \N__4964\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6131\,
            ce => \N__4209\,
            sr => \N__5816\
        );

    \fsm_ctrl_inst1.current_state_RNI2HR8_1_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4961\,
            lcout => \fsm_ctrl_inst1.current_state_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.bit_sequence_din_3_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3195\,
            in2 => \_gnd_net_\,
            in3 => \N__4591\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6136\,
            ce => \N__3326\,
            sr => \N__5820\
        );

    \fsm_ctrl_inst1.bit_sequence_din_5_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4595\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3279\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6136\,
            ce => \N__3326\,
            sr => \N__5820\
        );

    \fsm_ctrl_inst1.bit_sequence_din_10_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3381\,
            in2 => \_gnd_net_\,
            in3 => \N__4590\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6136\,
            ce => \N__3326\,
            sr => \N__5820\
        );

    \fsm_ctrl_inst1.bit_sequence_din_2_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4594\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3204\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6136\,
            ce => \N__3326\,
            sr => \N__5820\
        );

    \fsm_ctrl_inst1.bit_sequence_din_6_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3189\,
            in2 => \_gnd_net_\,
            in3 => \N__4593\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6136\,
            ce => \N__3326\,
            sr => \N__5820\
        );

    \fsm_ctrl_inst1.bit_sequence_din_4_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3285\,
            in2 => \_gnd_net_\,
            in3 => \N__4592\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6136\,
            ce => \N__3326\,
            sr => \N__5820\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_56_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3261\,
            in2 => \_gnd_net_\,
            in3 => \N__5038\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6120\,
            ce => \N__4199\,
            sr => \N__5805\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_60_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5039\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3267\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6120\,
            ce => \N__4199\,
            sr => \N__5805\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_55_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3411\,
            in2 => \_gnd_net_\,
            in3 => \N__5037\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6120\,
            ce => \N__4199\,
            sr => \N__5805\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_8_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4970\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3255\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6125\,
            ce => \N__4204\,
            sr => \N__5808\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_10_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3243\,
            in2 => \_gnd_net_\,
            in3 => \N__4967\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6125\,
            ce => \N__4204\,
            sr => \N__5808\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_9_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3249\,
            in2 => \_gnd_net_\,
            in3 => \N__4971\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6125\,
            ce => \N__4204\,
            sr => \N__5808\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_11_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4968\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3237\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6125\,
            ce => \N__4204\,
            sr => \N__5808\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_83_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3444\,
            in2 => \_gnd_net_\,
            in3 => \N__4969\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6125\,
            ce => \N__4204\,
            sr => \N__5808\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_42_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__3495\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4965\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6128\,
            ce => \N__4206\,
            sr => \N__5812\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_43_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3303\,
            in2 => \_gnd_net_\,
            in3 => \N__4966\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6128\,
            ce => \N__4206\,
            sr => \N__5812\
        );

    \fsm_ctrl_inst1.counter_idle_cry_c_0_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4042\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_20_0_\,
            carryout => \fsm_ctrl_inst1.counter_idle_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_RNO_0_1_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4116\,
            in2 => \_gnd_net_\,
            in3 => \N__3297\,
            lcout => \fsm_ctrl_inst1.counter_idle_s_1\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_idle_cry_0\,
            carryout => \fsm_ctrl_inst1.counter_idle_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_RNO_0_2_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3966\,
            in2 => \_gnd_net_\,
            in3 => \N__3294\,
            lcout => \fsm_ctrl_inst1.counter_idle_s_2\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_idle_cry_1\,
            carryout => \fsm_ctrl_inst1.counter_idle_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_RNO_0_3_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4075\,
            in2 => \_gnd_net_\,
            in3 => \N__3291\,
            lcout => \fsm_ctrl_inst1.counter_idle_s_3\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_idle_cry_2\,
            carryout => \fsm_ctrl_inst1.counter_idle_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_RNO_0_4_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4010\,
            in2 => \_gnd_net_\,
            in3 => \N__3288\,
            lcout => \fsm_ctrl_inst1.counter_idle_s_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_RNO_2_1_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__4012\,
            in1 => \N__3972\,
            in2 => \N__4960\,
            in3 => \N__4543\,
            lcout => \fsm_ctrl_inst1.g0_0_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_din_0_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4267\,
            in2 => \_gnd_net_\,
            in3 => \N__4544\,
            lcout => \fsm_ctrl_inst1.counter_dinZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6137\,
            ce => 'H',
            sr => \N__5821\
        );

    \fsm_ctrl_inst1.counter_idle_RNO_1_1_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4084\,
            in2 => \_gnd_net_\,
            in3 => \N__4119\,
            lcout => \fsm_ctrl_inst1.g0_0_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.bit_sequence_din_9_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4548\,
            in2 => \_gnd_net_\,
            in3 => \N__3363\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6141\,
            ce => \N__3327\,
            sr => \N__5826\
        );

    \fsm_ctrl_inst1.bit_sequence_din_12_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4549\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3345\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6141\,
            ce => \N__3327\,
            sr => \N__5826\
        );

    \fsm_ctrl_inst1.bit_sequence_din_7_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4547\,
            in2 => \_gnd_net_\,
            in3 => \N__3375\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6141\,
            ce => \N__3327\,
            sr => \N__5826\
        );

    \fsm_ctrl_inst1.bit_sequence_din_8_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4552\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3369\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6141\,
            ce => \N__3327\,
            sr => \N__5826\
        );

    \fsm_ctrl_inst1.bit_sequence_din_13_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4546\,
            in2 => \_gnd_net_\,
            in3 => \N__3357\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6141\,
            ce => \N__3327\,
            sr => \N__5826\
        );

    \fsm_ctrl_inst1.bit_sequence_din_15_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4551\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3333\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6141\,
            ce => \N__3327\,
            sr => \N__5826\
        );

    \fsm_ctrl_inst1.bit_sequence_din_11_LC_3_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4545\,
            in2 => \_gnd_net_\,
            in3 => \N__3351\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6141\,
            ce => \N__3327\,
            sr => \N__5826\
        );

    \fsm_ctrl_inst1.bit_sequence_din_14_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4550\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3339\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6141\,
            ce => \N__3327\,
            sr => \N__5826\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_75_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5022\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3690\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6132\,
            ce => \N__4210\,
            sr => \N__5809\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_76_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3438\,
            in2 => \_gnd_net_\,
            in3 => \N__5023\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6132\,
            ce => \N__4210\,
            sr => \N__5809\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_77_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__5024\,
            in1 => \N__3432\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6132\,
            ce => \N__4210\,
            sr => \N__5809\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_78_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5011\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3426\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6129\,
            ce => \N__4207\,
            sr => \N__5803\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_12_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3420\,
            in2 => \_gnd_net_\,
            in3 => \N__5010\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6129\,
            ce => \N__4207\,
            sr => \N__5803\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_54_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3462\,
            in2 => \_gnd_net_\,
            in3 => \N__5000\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6123\,
            ce => \N__4202\,
            sr => \N__5810\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_62_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5002\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3399\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6123\,
            ce => \N__4202\,
            sr => \N__5810\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_80_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5004\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3387\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6123\,
            ce => \N__4202\,
            sr => \N__5810\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_61_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3405\,
            in2 => \_gnd_net_\,
            in3 => \N__5001\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6123\,
            ce => \N__4202\,
            sr => \N__5810\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_79_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5003\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3393\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6123\,
            ce => \N__4202\,
            sr => \N__5810\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_4_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3537\,
            in2 => \_gnd_net_\,
            in3 => \N__4988\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6130\,
            ce => \N__4208\,
            sr => \N__5813\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_81_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4991\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3483\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6130\,
            ce => \N__4208\,
            sr => \N__5813\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_37_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3852\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4985\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6130\,
            ce => \N__4208\,
            sr => \N__5813\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_5_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4990\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3477\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6130\,
            ce => \N__4208\,
            sr => \N__5813\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_48_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3813\,
            in2 => \_gnd_net_\,
            in3 => \N__4987\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6130\,
            ce => \N__4208\,
            sr => \N__5813\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_53_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4989\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3789\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6130\,
            ce => \N__4208\,
            sr => \N__5813\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_38_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3456\,
            in2 => \_gnd_net_\,
            in3 => \N__4986\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6130\,
            ce => \N__4208\,
            sr => \N__5813\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_82_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4992\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3450\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6130\,
            ce => \N__4208\,
            sr => \N__5813\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_40_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4858\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3513\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6133\,
            ce => \N__4211\,
            sr => \N__5817\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_1_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3507\,
            in2 => \_gnd_net_\,
            in3 => \N__4854\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6133\,
            ce => \N__4211\,
            sr => \N__5817\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_3_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4857\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3525\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6133\,
            ce => \N__4211\,
            sr => \N__5817\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_2_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3531\,
            in2 => \_gnd_net_\,
            in3 => \N__4855\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6133\,
            ce => \N__4211\,
            sr => \N__5817\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_39_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4856\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3519\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6133\,
            ce => \N__4211\,
            sr => \N__5817\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_0_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4853\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6133\,
            ce => \N__4211\,
            sr => \N__5817\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_41_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4859\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3501\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6133\,
            ce => \N__4211\,
            sr => \N__5817\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_44_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3489\,
            in2 => \_gnd_net_\,
            in3 => \N__4860\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6133\,
            ce => \N__4211\,
            sr => \N__5817\
        );

    \fsm_ctrl_inst1.counter_idle_RNO_2_2_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__4011\,
            in1 => \N__4542\,
            in2 => \N__4808\,
            in3 => \N__3969\,
            lcout => \fsm_ctrl_inst1.g0_0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_RNO_1_2_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4077\,
            in2 => \_gnd_net_\,
            in3 => \N__4120\,
            lcout => \fsm_ctrl_inst1.g0_0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_RNO_1_3_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__4121\,
            in1 => \_gnd_net_\,
            in2 => \N__4085\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.g0_0_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_3_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__4020\,
            in1 => \N__3636\,
            in2 => \N__3579\,
            in3 => \N__3576\,
            lcout => \fsm_ctrl_inst1.counter_idleZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6138\,
            ce => 'H',
            sr => \N__5822\
        );

    \fsm_ctrl_inst1.counter_idle_RNO_1_4_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__4122\,
            in1 => \_gnd_net_\,
            in2 => \N__4086\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.g0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_4_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__3936\,
            in1 => \N__3637\,
            in2 => \N__3570\,
            in3 => \N__3567\,
            lcout => \fsm_ctrl_inst1.counter_idleZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6138\,
            ce => 'H',
            sr => \N__5822\
        );

    \fsm_ctrl_inst1.current_state_RNI31NH_0_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__4690\,
            in1 => \N__4541\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_ctrl_inst1.current_state_20_d_i\,
            ltout => \fsm_ctrl_inst1.current_state_20_d_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_2_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000111110001000"
        )
    port map (
            in0 => \N__3561\,
            in1 => \N__3555\,
            in2 => \N__3549\,
            in3 => \N__3546\,
            lcout => \fsm_ctrl_inst1.counter_idleZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6138\,
            ce => 'H',
            sr => \N__5822\
        );

    \fsm_ctrl_inst1.current_state_RNO_0_0_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3968\,
            in2 => \_gnd_net_\,
            in3 => \N__4026\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.N_93_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.current_state_0_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__4852\,
            in1 => \N__3924\,
            in2 => \N__3540\,
            in3 => \N__4584\,
            lcout => fsm_ctrl_inst1_current_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6142\,
            ce => 'H',
            sr => \N__5827\
        );

    \fsm_ctrl_inst1.counter_idle_RNO_1_0_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4076\,
            in1 => \N__3967\,
            in2 => \N__4014\,
            in3 => \N__4118\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.counter_idle_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_RNO_0_0_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4694\,
            in2 => \N__3666\,
            in3 => \N__4583\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.counter_idlee_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_0_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000100000100"
        )
    port map (
            in0 => \N__3639\,
            in1 => \N__3600\,
            in2 => \N__3663\,
            in3 => \N__4044\,
            lcout => \fsm_ctrl_inst1.counter_idleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6142\,
            ce => 'H',
            sr => \N__5827\
        );

    \fsm_ctrl_inst1.counter_idle_1_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__3660\,
            in1 => \N__3654\,
            in2 => \N__3648\,
            in3 => \N__3638\,
            lcout => \fsm_ctrl_inst1.counter_idleZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6142\,
            ce => 'H',
            sr => \N__5827\
        );

    \fsm_ctrl_inst1.MOSI_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__3621\,
            in1 => \N__4553\,
            in2 => \N__3615\,
            in3 => \N__4807\,
            lcout => \MOSI\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6144\,
            ce => 'H',
            sr => \N__5828\
        );

    \CONSTANT_ONE_LUT4_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_67_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5052\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3720\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6145\,
            ce => \N__4217\,
            sr => \N__5823\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_68_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3591\,
            in2 => \_gnd_net_\,
            in3 => \N__5053\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6145\,
            ce => \N__4217\,
            sr => \N__5823\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_65_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5050\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3585\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6145\,
            ce => \N__4217\,
            sr => \N__5823\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_64_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3753\,
            in2 => \_gnd_net_\,
            in3 => \N__5049\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6145\,
            ce => \N__4217\,
            sr => \N__5823\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_66_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5051\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3726\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6145\,
            ce => \N__4217\,
            sr => \N__5823\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_69_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3714\,
            in2 => \_gnd_net_\,
            in3 => \N__5045\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6143\,
            ce => \N__4216\,
            sr => \N__5818\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_70_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3708\,
            in2 => \_gnd_net_\,
            in3 => \N__5046\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6143\,
            ce => \N__4216\,
            sr => \N__5818\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_71_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5047\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3702\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6143\,
            ce => \N__4216\,
            sr => \N__5818\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_73_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3678\,
            in2 => \_gnd_net_\,
            in3 => \N__5008\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6139\,
            ce => \N__4214\,
            sr => \N__5814\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_74_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5009\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3696\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6139\,
            ce => \N__4214\,
            sr => \N__5814\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_19_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3672\,
            in2 => \_gnd_net_\,
            in3 => \N__5006\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6139\,
            ce => \N__4214\,
            sr => \N__5814\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_72_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5007\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3684\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6139\,
            ce => \N__4214\,
            sr => \N__5814\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_18_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3783\,
            in2 => \_gnd_net_\,
            in3 => \N__5005\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6139\,
            ce => \N__4214\,
            sr => \N__5814\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_14_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3831\,
            in2 => \_gnd_net_\,
            in3 => \N__4993\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6134\,
            ce => \N__4212\,
            sr => \N__5806\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_17_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4996\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3777\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6134\,
            ce => \N__4212\,
            sr => \N__5806\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_16_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3765\,
            in2 => \_gnd_net_\,
            in3 => \N__4995\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6134\,
            ce => \N__4212\,
            sr => \N__5806\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_21_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4997\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4227\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6134\,
            ce => \N__4212\,
            sr => \N__5806\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_15_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__4994\,
            in1 => \N__3771\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6134\,
            ce => \N__4212\,
            sr => \N__5806\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_63_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3759\,
            in2 => \_gnd_net_\,
            in3 => \N__4999\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6134\,
            ce => \N__4212\,
            sr => \N__5806\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_22_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4998\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3744\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6134\,
            ce => \N__4212\,
            sr => \N__5806\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_27_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3846\,
            in2 => \_gnd_net_\,
            in3 => \N__4953\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6126\,
            ce => \N__4205\,
            sr => \N__5815\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_23_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4951\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3738\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6126\,
            ce => \N__4205\,
            sr => \N__5815\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_49_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3732\,
            in2 => \_gnd_net_\,
            in3 => \N__4954\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6126\,
            ce => \N__4205\,
            sr => \N__5815\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_26_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4952\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3807\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6126\,
            ce => \N__4205\,
            sr => \N__5815\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_13_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3840\,
            in2 => \_gnd_net_\,
            in3 => \N__4950\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6126\,
            ce => \N__4205\,
            sr => \N__5815\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_50_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3825\,
            in2 => \_gnd_net_\,
            in3 => \N__4955\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6126\,
            ce => \N__4205\,
            sr => \N__5815\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_51_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4956\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3819\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6126\,
            ce => \N__4205\,
            sr => \N__5815\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_47_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4948\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3900\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6135\,
            ce => \N__4213\,
            sr => \N__5819\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_25_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3912\,
            in2 => \_gnd_net_\,
            in3 => \N__4943\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6135\,
            ce => \N__4213\,
            sr => \N__5819\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_45_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4946\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3801\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6135\,
            ce => \N__4213\,
            sr => \N__5819\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_29_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3888\,
            in2 => \_gnd_net_\,
            in3 => \N__4945\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6135\,
            ce => \N__4213\,
            sr => \N__5819\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_52_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4949\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3795\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6135\,
            ce => \N__4213\,
            sr => \N__5819\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_24_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3918\,
            in2 => \_gnd_net_\,
            in3 => \N__4942\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6135\,
            ce => \N__4213\,
            sr => \N__5819\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_46_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4947\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3906\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6135\,
            ce => \N__4213\,
            sr => \N__5819\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_28_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3894\,
            in2 => \_gnd_net_\,
            in3 => \N__4944\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6135\,
            ce => \N__4213\,
            sr => \N__5819\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_33_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4128\,
            in2 => \_gnd_net_\,
            in3 => \N__4864\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6140\,
            ce => \N__4215\,
            sr => \N__5824\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_34_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4865\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3882\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6140\,
            ce => \N__4215\,
            sr => \N__5824\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_30_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3876\,
            in2 => \_gnd_net_\,
            in3 => \N__4861\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6140\,
            ce => \N__4215\,
            sr => \N__5824\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_35_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4866\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3870\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6140\,
            ce => \N__4215\,
            sr => \N__5824\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_31_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4862\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3864\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6140\,
            ce => \N__4215\,
            sr => \N__5824\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_36_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3858\,
            in2 => \_gnd_net_\,
            in3 => \N__4867\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6140\,
            ce => \N__4215\,
            sr => \N__5824\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_32_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4863\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4134\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6140\,
            ce => \N__4215\,
            sr => \N__5824\
        );

    \fsm_ctrl_inst1.current_state_RNO_2_0_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4117\,
            in1 => \N__4074\,
            in2 => \N__4013\,
            in3 => \N__4043\,
            lcout => \fsm_ctrl_inst1.current_state_RNO_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_RNO_2_3_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__4005\,
            in1 => \N__3970\,
            in2 => \N__4809\,
            in3 => \N__4508\,
            lcout => \fsm_ctrl_inst1.g0_0_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst1.STATSR_cnv_x0_0_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5093\,
            in1 => \N__4439\,
            in2 => \N__5076\,
            in3 => \N__4507\,
            lcout => \config_register_latched_dec_inst1.STATSR_cnv_x0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_RNO_2_4_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__4006\,
            in1 => \N__3971\,
            in2 => \N__4810\,
            in3 => \N__4509\,
            lcout => \fsm_ctrl_inst1.g0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_din_RNO_0_3_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__4327\,
            in1 => \N__4272\,
            in2 => \N__4313\,
            in3 => \N__4287\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.counter_din_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_din_3_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__4567\,
            in1 => \_gnd_net_\,
            in2 => \N__3930\,
            in3 => \_gnd_net_\,
            lcout => \fsm_ctrl_inst1.counter_dinZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6146\,
            ce => 'H',
            sr => \N__5829\
        );

    \fsm_ctrl_inst1.current_state_RNO_3_0_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4326\,
            in1 => \N__4565\,
            in2 => \N__4312\,
            in3 => \N__4286\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.current_state_RNO_3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.current_state_RNO_1_0_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3927\,
            in3 => \N__4268\,
            lcout => \fsm_ctrl_inst1.current_state_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_din_1_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__4269\,
            in1 => \N__4569\,
            in2 => \_gnd_net_\,
            in3 => \N__4288\,
            lcout => \fsm_ctrl_inst1.counter_dinZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6146\,
            ce => 'H',
            sr => \N__5829\
        );

    \fsm_ctrl_inst1.counter_din_2_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010101010000000"
        )
    port map (
            in0 => \N__4568\,
            in1 => \N__4270\,
            in2 => \N__4293\,
            in3 => \N__4329\,
            lcout => \fsm_ctrl_inst1.counter_dinZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6146\,
            ce => 'H',
            sr => \N__5829\
        );

    \fsm_ctrl_inst1.current_state_RNO_0_1_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__4328\,
            in1 => \_gnd_net_\,
            in2 => \N__4314\,
            in3 => \N__4566\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.o2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.current_state_1_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__4292\,
            in1 => \N__4271\,
            in2 => \N__4242\,
            in3 => \N__4806\,
            lcout => fsm_ctrl_inst1_current_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6146\,
            ce => 'H',
            sr => \N__5829\
        );

    \config_register_latched_dec_inst1.STATSR_0_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4418\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6150\,
            ce => \N__5976\,
            sr => \N__5832\
        );

    \config_register_latched_dec_inst1.STATSR_1_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4239\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6153\,
            ce => \N__5975\,
            sr => \N__5835\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_20_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4233\,
            in2 => \_gnd_net_\,
            in3 => \N__5048\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6147\,
            ce => \N__4218\,
            sr => \N__5825\
        );

    \config_register_latched_dec_inst1.DYNSR_RNIQ2U9_15_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4368\,
            in1 => \N__5202\,
            in2 => \_gnd_net_\,
            in3 => \N__4446\,
            lcout => \SDO_signal_out_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst1.DYNSR_12_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4344\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6148\,
            ce => \N__5145\,
            sr => \N__5830\
        );

    \config_register_latched_dec_inst1.DYNSR_14_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4356\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6148\,
            ce => \N__5145\,
            sr => \N__5830\
        );

    \config_register_latched_dec_inst1.DYNSR_10_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5193\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6148\,
            ce => \N__5145\,
            sr => \N__5830\
        );

    \config_register_latched_dec_inst1.DYNSR_15_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4374\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6148\,
            ce => \N__5145\,
            sr => \N__5830\
        );

    \config_register_latched_dec_inst1.DYNSR_13_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4362\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6148\,
            ce => \N__5145\,
            sr => \N__5830\
        );

    \config_register_latched_dec_inst1.DYNSR_11_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4350\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6148\,
            ce => \N__5145\,
            sr => \N__5830\
        );

    \config_register_latched_dec_inst1.DYNSR_cnv_x0_0_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__4554\,
            in1 => \N__5075\,
            in2 => \N__5115\,
            in3 => \N__4442\,
            lcout => OPEN,
            ltout => \config_register_latched_dec_inst1.DYNSR_cnv_x0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst1.DYNSR_cnv_ns_0_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4335\,
            in2 => \N__4338\,
            in3 => \N__4688\,
            lcout => \config_register_latched_dec_inst1.DYNSR_cnv_nsZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst1.DYNSR_cnv_x1_0_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5112\,
            in1 => \N__5073\,
            in2 => \_gnd_net_\,
            in3 => \N__4440\,
            lcout => \config_register_latched_dec_inst1.DYNSR_cnv_x1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.SCLK_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__5114\,
            in1 => \N__4689\,
            in2 => \_gnd_net_\,
            in3 => \N__4556\,
            lcout => \fsm_ctrl_inst1_SCLK_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6149\,
            ce => 'H',
            sr => \N__5831\
        );

    \config_register_latched_dec_inst1.STATSR_cnv_x1_0_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__5113\,
            in1 => \N__4441\,
            in2 => \_gnd_net_\,
            in3 => \N__5074\,
            lcout => OPEN,
            ltout => \config_register_latched_dec_inst1.STATSR_cnv_x1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst1.STATSR_cnv_ns_0_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4687\,
            in2 => \N__4617\,
            in3 => \N__4614\,
            lcout => \STATSR_cnv_ns_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.SEL_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4555\,
            lcout => \SEL_REG\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6149\,
            ce => 'H',
            sr => \N__5831\
        );

    \config_register_latched_dec_inst1.DYNSR_2_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4398\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6151\,
            ce => \N__5153\,
            sr => \N__5833\
        );

    \config_register_latched_dec_inst1.DYNSR_0_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4419\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6151\,
            ce => \N__5153\,
            sr => \N__5833\
        );

    \config_register_latched_dec_inst1.DYNSR_1_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4404\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6151\,
            ce => \N__5153\,
            sr => \N__5833\
        );

    \config_register_latched_dec_inst1.DYNSR_3_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4392\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6151\,
            ce => \N__5153\,
            sr => \N__5833\
        );

    \config_register_latched_dec_inst1.DYNSR_4_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4386\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6151\,
            ce => \N__5153\,
            sr => \N__5833\
        );

    \config_register_latched_dec_inst1.STATSR_2_LC_6_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4380\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6155\,
            ce => \N__5974\,
            sr => \N__5837\
        );

    \config_register_latched_dec_inst1.STATSR_3_LC_6_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5214\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6155\,
            ce => \N__5974\,
            sr => \N__5837\
        );

    \config_register_latched_dec_inst1.STATSR_4_LC_6_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5208\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6155\,
            ce => \N__5974\,
            sr => \N__5837\
        );

    \config_register_latched_dec_inst1.STATSR_87_LC_6_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5262\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6156\,
            ce => \N__5972\,
            sr => \N__5838\
        );

    \config_register_latched_dec_inst1.DYNSR_9_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5175\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6152\,
            ce => \N__5157\,
            sr => \N__5834\
        );

    \config_register_latched_dec_inst1.DYNSR_6_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5163\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6152\,
            ce => \N__5157\,
            sr => \N__5834\
        );

    \config_register_latched_dec_inst1.DYNSR_7_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5187\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6152\,
            ce => \N__5157\,
            sr => \N__5834\
        );

    \config_register_latched_dec_inst1.DYNSR_8_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5181\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6152\,
            ce => \N__5157\,
            sr => \N__5834\
        );

    \config_register_latched_dec_inst1.DYNSR_5_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5169\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6154\,
            ce => \N__5152\,
            sr => \N__5836\
        );

    \config_register_latched_dec_inst1.STATSR_6_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5268\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6157\,
            ce => \N__5973\,
            sr => \N__5839\
        );

    \config_register_latched_dec_inst1.STATSR_5_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5274\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6157\,
            ce => \N__5973\,
            sr => \N__5839\
        );

    \config_register_latched_dec_inst1.STATSR_86_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5229\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6158\,
            ce => \N__5971\,
            sr => \N__5840\
        );

    \config_register_latched_dec_inst1.STATSR_8_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5247\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6159\,
            ce => \N__5970\,
            sr => \N__5841\
        );

    \config_register_latched_dec_inst1.STATSR_7_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5256\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6159\,
            ce => \N__5970\,
            sr => \N__5841\
        );

    \config_register_latched_dec_inst1.STATSR_84_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5316\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6160\,
            ce => \N__5969\,
            sr => \N__5842\
        );

    \config_register_latched_dec_inst1.STATSR_9_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5241\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6160\,
            ce => \N__5969\,
            sr => \N__5842\
        );

    \config_register_latched_dec_inst1.STATSR_85_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5235\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6160\,
            ce => \N__5969\,
            sr => \N__5842\
        );

    \config_register_latched_dec_inst1.STATSR_12_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5322\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6161\,
            ce => \N__5968\,
            sr => \N__5843\
        );

    \config_register_latched_dec_inst1.STATSR_10_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5220\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6161\,
            ce => \N__5968\,
            sr => \N__5843\
        );

    \config_register_latched_dec_inst1.STATSR_11_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5328\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6161\,
            ce => \N__5968\,
            sr => \N__5843\
        );

    \config_register_latched_dec_inst1.STATSR_83_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5298\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6162\,
            ce => \N__5966\,
            sr => \N__5844\
        );

    \config_register_latched_dec_inst1.STATSR_13_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5310\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6163\,
            ce => \N__5967\,
            sr => \N__5845\
        );

    \config_register_latched_dec_inst1.STATSR_81_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5286\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6164\,
            ce => \N__5964\,
            sr => \N__5846\
        );

    \config_register_latched_dec_inst1.STATSR_82_LC_11_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5304\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6164\,
            ce => \N__5964\,
            sr => \N__5846\
        );

    \config_register_latched_dec_inst1.STATSR_14_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5292\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6165\,
            ce => \N__5965\,
            sr => \N__5847\
        );

    \config_register_latched_dec_inst1.STATSR_77_LC_12_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5364\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6167\,
            ce => \N__5961\,
            sr => \N__5849\
        );

    \config_register_latched_dec_inst1.STATSR_80_LC_12_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5280\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6167\,
            ce => \N__5961\,
            sr => \N__5849\
        );

    \config_register_latched_dec_inst1.STATSR_79_LC_12_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5382\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6167\,
            ce => \N__5961\,
            sr => \N__5849\
        );

    \config_register_latched_dec_inst1.STATSR_78_LC_12_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5388\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6167\,
            ce => \N__5961\,
            sr => \N__5849\
        );

    \config_register_latched_dec_inst1.STATSR_15_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5376\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6166\,
            ce => \N__5963\,
            sr => \N__5848\
        );

    \config_register_latched_dec_inst1.STATSR_75_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5358\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6169\,
            ce => \N__5959\,
            sr => \N__5851\
        );

    \config_register_latched_dec_inst1.STATSR_76_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5370\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6169\,
            ce => \N__5959\,
            sr => \N__5851\
        );

    \config_register_latched_dec_inst1.STATSR_74_LC_13_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5340\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6171\,
            ce => \N__5957\,
            sr => \N__5853\
        );

    \config_register_latched_dec_inst1.STATSR_16_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5352\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6168\,
            ce => \N__5962\,
            sr => \N__5850\
        );

    \config_register_latched_dec_inst1.STATSR_17_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5346\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6170\,
            ce => \N__5960\,
            sr => \N__5852\
        );

    \config_register_latched_dec_inst1.STATSR_73_LC_14_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5424\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6173\,
            ce => \N__5956\,
            sr => \N__5855\
        );

    \config_register_latched_dec_inst1.STATSR_18_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5334\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6172\,
            ce => \N__5958\,
            sr => \N__5854\
        );

    \config_register_latched_dec_inst1.STATSR_19_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5436\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6172\,
            ce => \N__5958\,
            sr => \N__5854\
        );

    \config_register_latched_dec_inst1.STATSR_71_LC_15_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5418\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6174\,
            ce => \N__5953\,
            sr => \N__5856\
        );

    \config_register_latched_dec_inst1.STATSR_72_LC_15_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5430\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6174\,
            ce => \N__5953\,
            sr => \N__5856\
        );

    \config_register_latched_dec_inst1.STATSR_70_LC_15_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5406\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6176\,
            ce => \N__5950\,
            sr => \N__5858\
        );

    \config_register_latched_dec_inst1.STATSR_68_LC_15_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5400\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6176\,
            ce => \N__5950\,
            sr => \N__5858\
        );

    \config_register_latched_dec_inst1.STATSR_69_LC_15_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5412\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6176\,
            ce => \N__5950\,
            sr => \N__5858\
        );

    \config_register_latched_dec_inst1.STATSR_67_LC_15_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5394\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6176\,
            ce => \N__5950\,
            sr => \N__5858\
        );

    \config_register_latched_dec_inst1.STATSR_66_LC_15_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5442\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6179\,
            ce => \N__5948\,
            sr => \N__5861\
        );

    \config_register_latched_dec_inst1.STATSR_21_LC_16_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5490\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6175\,
            ce => \N__5954\,
            sr => \N__5857\
        );

    \config_register_latched_dec_inst1.STATSR_20_LC_16_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5496\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6175\,
            ce => \N__5954\,
            sr => \N__5857\
        );

    \config_register_latched_dec_inst1.STATSR_41_LC_16_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5478\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6175\,
            ce => \N__5954\,
            sr => \N__5857\
        );

    \config_register_latched_dec_inst1.STATSR_42_LC_16_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5484\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6175\,
            ce => \N__5954\,
            sr => \N__5857\
        );

    \config_register_latched_dec_inst1.STATSR_40_LC_16_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5526\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6175\,
            ce => \N__5954\,
            sr => \N__5857\
        );

    \config_register_latched_dec_inst1.STATSR_44_LC_16_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5466\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6177\,
            ce => \N__5951\,
            sr => \N__5859\
        );

    \config_register_latched_dec_inst1.STATSR_43_LC_16_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5472\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6177\,
            ce => \N__5951\,
            sr => \N__5859\
        );

    \config_register_latched_dec_inst1.STATSR_45_LC_16_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5460\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6177\,
            ce => \N__5951\,
            sr => \N__5859\
        );

    \config_register_latched_dec_inst1.STATSR_46_LC_16_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5454\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6177\,
            ce => \N__5951\,
            sr => \N__5859\
        );

    \config_register_latched_dec_inst1.STATSR_22_LC_16_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5448\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6177\,
            ce => \N__5951\,
            sr => \N__5859\
        );

    \config_register_latched_dec_inst1.STATSR_65_LC_16_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5568\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6182\,
            ce => \N__5945\,
            sr => \N__5864\
        );

    \config_register_latched_dec_inst1.STATSR_36_LC_17_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5544\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6178\,
            ce => \N__5949\,
            sr => \N__5860\
        );

    \config_register_latched_dec_inst1.STATSR_37_LC_17_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5550\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6178\,
            ce => \N__5949\,
            sr => \N__5860\
        );

    \config_register_latched_dec_inst1.STATSR_35_LC_17_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5640\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6178\,
            ce => \N__5949\,
            sr => \N__5860\
        );

    \config_register_latched_dec_inst1.STATSR_38_LC_17_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5538\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6178\,
            ce => \N__5949\,
            sr => \N__5860\
        );

    \config_register_latched_dec_inst1.STATSR_39_LC_17_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5532\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6178\,
            ce => \N__5949\,
            sr => \N__5860\
        );

    \config_register_latched_dec_inst1.STATSR_47_LC_17_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5520\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6180\,
            ce => \N__5947\,
            sr => \N__5862\
        );

    \config_register_latched_dec_inst1.STATSR_48_LC_17_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5514\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6180\,
            ce => \N__5947\,
            sr => \N__5862\
        );

    \config_register_latched_dec_inst1.STATSR_23_LC_17_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5508\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6180\,
            ce => \N__5947\,
            sr => \N__5862\
        );

    \config_register_latched_dec_inst1.STATSR_49_LC_17_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5502\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6180\,
            ce => \N__5947\,
            sr => \N__5862\
        );

    \config_register_latched_dec_inst1.STATSR_24_LC_17_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5598\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6180\,
            ce => \N__5947\,
            sr => \N__5862\
        );

    \config_register_latched_dec_inst1.STATSR_50_LC_17_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5592\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6183\,
            ce => \N__5944\,
            sr => \N__5865\
        );

    \config_register_latched_dec_inst1.STATSR_52_LC_17_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5574\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6183\,
            ce => \N__5944\,
            sr => \N__5865\
        );

    \config_register_latched_dec_inst1.STATSR_53_LC_17_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5586\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6183\,
            ce => \N__5944\,
            sr => \N__5865\
        );

    \config_register_latched_dec_inst1.STATSR_51_LC_17_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5580\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6183\,
            ce => \N__5944\,
            sr => \N__5865\
        );

    \config_register_latched_dec_inst1.STATSR_64_LC_17_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5562\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6185\,
            ce => \N__5943\,
            sr => \N__5867\
        );

    \config_register_latched_dec_inst1.STATSR_63_LC_17_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5652\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6185\,
            ce => \N__5943\,
            sr => \N__5867\
        );

    \config_register_latched_dec_inst1.STATSR_61_LC_17_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6228\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6185\,
            ce => \N__5943\,
            sr => \N__5867\
        );

    \config_register_latched_dec_inst1.STATSR_54_LC_17_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5556\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6185\,
            ce => \N__5943\,
            sr => \N__5867\
        );

    \config_register_latched_dec_inst1.STATSR_62_LC_17_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5658\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6185\,
            ce => \N__5943\,
            sr => \N__5867\
        );

    \config_register_latched_dec_inst1.STATSR_31_LC_18_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5646\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6181\,
            ce => \N__5955\,
            sr => \N__5863\
        );

    \config_register_latched_dec_inst1.STATSR_30_LC_18_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6234\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6181\,
            ce => \N__5955\,
            sr => \N__5863\
        );

    \config_register_latched_dec_inst1.STATSR_34_LC_18_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5622\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6181\,
            ce => \N__5955\,
            sr => \N__5863\
        );

    \config_register_latched_dec_inst1.STATSR_32_LC_18_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5634\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6181\,
            ce => \N__5955\,
            sr => \N__5863\
        );

    \config_register_latched_dec_inst1.STATSR_33_LC_18_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5628\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6181\,
            ce => \N__5955\,
            sr => \N__5863\
        );

    \config_register_latched_dec_inst1.STATSR_26_LC_18_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5604\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6184\,
            ce => \N__5952\,
            sr => \N__5866\
        );

    \config_register_latched_dec_inst1.STATSR_27_LC_18_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5616\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6184\,
            ce => \N__5952\,
            sr => \N__5866\
        );

    \config_register_latched_dec_inst1.STATSR_25_LC_18_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5610\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6184\,
            ce => \N__5952\,
            sr => \N__5866\
        );

    \config_register_latched_dec_inst1.STATSR_28_LC_18_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6246\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6184\,
            ce => \N__5952\,
            sr => \N__5866\
        );

    \config_register_latched_dec_inst1.STATSR_29_LC_18_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6240\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6184\,
            ce => \N__5952\,
            sr => \N__5866\
        );

    \config_register_latched_dec_inst1.STATSR_60_LC_18_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6216\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6186\,
            ce => \N__5946\,
            sr => \N__5868\
        );

    \config_register_latched_dec_inst1.STATSR_55_LC_18_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6222\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6186\,
            ce => \N__5946\,
            sr => \N__5868\
        );

    \config_register_latched_dec_inst1.STATSR_59_LC_18_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6204\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6186\,
            ce => \N__5946\,
            sr => \N__5868\
        );

    \config_register_latched_dec_inst1.STATSR_57_LC_18_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6192\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6186\,
            ce => \N__5946\,
            sr => \N__5868\
        );

    \config_register_latched_dec_inst1.STATSR_58_LC_18_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6210\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6186\,
            ce => \N__5946\,
            sr => \N__5868\
        );

    \config_register_latched_dec_inst1.STATSR_56_LC_18_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6198\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6186\,
            ce => \N__5946\,
            sr => \N__5868\
        );
end \INTERFACE\;
