-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 13 2025 09:52:51

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    signal_out : out std_logic;
    CLK : in std_logic;
    SELSTAT : in std_logic;
    SELDYN : in std_logic;
    RST_N : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__2717\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2705\ : std_logic;
signal \N__2704\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2688\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2607\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2586\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2583\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2578\ : std_logic;
signal \N__2577\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2566\ : std_logic;
signal \N__2565\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2538\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2535\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2533\ : std_logic;
signal \N__2532\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2530\ : std_logic;
signal \N__2529\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2527\ : std_logic;
signal \N__2526\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2476\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2446\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2395\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2385\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2380\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2377\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2374\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2368\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2365\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2361\ : std_logic;
signal \N__2358\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2328\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2326\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2323\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2296\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2273\ : std_logic;
signal \N__2270\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2263\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2260\ : std_logic;
signal \N__2259\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2257\ : std_logic;
signal \N__2256\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2254\ : std_logic;
signal \N__2253\ : std_logic;
signal \N__2252\ : std_logic;
signal \N__2251\ : std_logic;
signal \N__2250\ : std_logic;
signal \N__2249\ : std_logic;
signal \N__2248\ : std_logic;
signal \N__2213\ : std_logic;
signal \N__2210\ : std_logic;
signal \N__2207\ : std_logic;
signal \N__2206\ : std_logic;
signal \N__2205\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2203\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2200\ : std_logic;
signal \N__2199\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2197\ : std_logic;
signal \N__2196\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2194\ : std_logic;
signal \N__2165\ : std_logic;
signal \N__2162\ : std_logic;
signal \N__2159\ : std_logic;
signal \N__2158\ : std_logic;
signal \N__2157\ : std_logic;
signal \N__2156\ : std_logic;
signal \N__2155\ : std_logic;
signal \N__2154\ : std_logic;
signal \N__2153\ : std_logic;
signal \N__2152\ : std_logic;
signal \N__2151\ : std_logic;
signal \N__2150\ : std_logic;
signal \N__2149\ : std_logic;
signal \N__2148\ : std_logic;
signal \N__2147\ : std_logic;
signal \N__2146\ : std_logic;
signal \N__2145\ : std_logic;
signal \N__2144\ : std_logic;
signal \N__2143\ : std_logic;
signal \N__2108\ : std_logic;
signal \N__2105\ : std_logic;
signal \N__2102\ : std_logic;
signal \N__2099\ : std_logic;
signal \N__2096\ : std_logic;
signal \N__2093\ : std_logic;
signal \N__2090\ : std_logic;
signal \N__2087\ : std_logic;
signal \N__2084\ : std_logic;
signal \N__2081\ : std_logic;
signal \N__2078\ : std_logic;
signal \N__2075\ : std_logic;
signal \N__2072\ : std_logic;
signal \N__2069\ : std_logic;
signal \N__2066\ : std_logic;
signal \N__2063\ : std_logic;
signal \N__2060\ : std_logic;
signal \N__2057\ : std_logic;
signal \N__2054\ : std_logic;
signal \N__2051\ : std_logic;
signal \N__2048\ : std_logic;
signal \N__2045\ : std_logic;
signal \N__2042\ : std_logic;
signal \N__2039\ : std_logic;
signal \N__2036\ : std_logic;
signal \N__2033\ : std_logic;
signal \N__2030\ : std_logic;
signal \N__2027\ : std_logic;
signal \N__2024\ : std_logic;
signal \N__2021\ : std_logic;
signal \N__2018\ : std_logic;
signal \N__2015\ : std_logic;
signal \N__2012\ : std_logic;
signal \N__2009\ : std_logic;
signal \N__2006\ : std_logic;
signal \N__2003\ : std_logic;
signal \N__2000\ : std_logic;
signal \N__1997\ : std_logic;
signal \N__1994\ : std_logic;
signal \N__1991\ : std_logic;
signal \N__1988\ : std_logic;
signal \N__1985\ : std_logic;
signal \N__1982\ : std_logic;
signal \N__1979\ : std_logic;
signal \N__1976\ : std_logic;
signal \N__1973\ : std_logic;
signal \N__1970\ : std_logic;
signal \N__1967\ : std_logic;
signal \N__1964\ : std_logic;
signal \N__1961\ : std_logic;
signal \N__1958\ : std_logic;
signal \N__1955\ : std_logic;
signal \N__1952\ : std_logic;
signal \N__1949\ : std_logic;
signal \N__1946\ : std_logic;
signal \N__1943\ : std_logic;
signal \N__1940\ : std_logic;
signal \N__1937\ : std_logic;
signal \N__1934\ : std_logic;
signal \N__1931\ : std_logic;
signal \N__1928\ : std_logic;
signal \N__1925\ : std_logic;
signal \N__1922\ : std_logic;
signal \N__1919\ : std_logic;
signal \N__1916\ : std_logic;
signal \N__1913\ : std_logic;
signal \N__1910\ : std_logic;
signal \N__1907\ : std_logic;
signal \N__1904\ : std_logic;
signal \N__1901\ : std_logic;
signal \N__1898\ : std_logic;
signal \N__1895\ : std_logic;
signal \N__1892\ : std_logic;
signal \N__1889\ : std_logic;
signal \N__1886\ : std_logic;
signal \N__1883\ : std_logic;
signal \N__1880\ : std_logic;
signal \N__1877\ : std_logic;
signal \N__1874\ : std_logic;
signal \N__1871\ : std_logic;
signal \N__1868\ : std_logic;
signal \N__1865\ : std_logic;
signal \N__1862\ : std_logic;
signal \N__1859\ : std_logic;
signal \N__1856\ : std_logic;
signal \N__1853\ : std_logic;
signal \N__1850\ : std_logic;
signal \N__1847\ : std_logic;
signal \N__1844\ : std_logic;
signal \N__1841\ : std_logic;
signal \N__1838\ : std_logic;
signal \N__1835\ : std_logic;
signal \N__1832\ : std_logic;
signal \N__1829\ : std_logic;
signal \N__1826\ : std_logic;
signal \N__1823\ : std_logic;
signal \N__1820\ : std_logic;
signal \N__1817\ : std_logic;
signal \N__1814\ : std_logic;
signal \N__1811\ : std_logic;
signal \N__1808\ : std_logic;
signal \N__1805\ : std_logic;
signal \N__1802\ : std_logic;
signal \N__1799\ : std_logic;
signal \N__1796\ : std_logic;
signal \N__1793\ : std_logic;
signal \N__1790\ : std_logic;
signal \N__1789\ : std_logic;
signal \N__1788\ : std_logic;
signal \N__1787\ : std_logic;
signal \N__1786\ : std_logic;
signal \N__1785\ : std_logic;
signal \N__1784\ : std_logic;
signal \N__1783\ : std_logic;
signal \N__1782\ : std_logic;
signal \N__1781\ : std_logic;
signal \N__1780\ : std_logic;
signal \N__1779\ : std_logic;
signal \N__1778\ : std_logic;
signal \N__1777\ : std_logic;
signal \N__1776\ : std_logic;
signal \N__1775\ : std_logic;
signal \N__1774\ : std_logic;
signal \N__1773\ : std_logic;
signal \N__1772\ : std_logic;
signal \N__1769\ : std_logic;
signal \N__1764\ : std_logic;
signal \N__1747\ : std_logic;
signal \N__1730\ : std_logic;
signal \N__1721\ : std_logic;
signal \N__1718\ : std_logic;
signal \N__1715\ : std_logic;
signal \N__1712\ : std_logic;
signal \N__1709\ : std_logic;
signal \N__1706\ : std_logic;
signal \N__1703\ : std_logic;
signal \N__1700\ : std_logic;
signal \N__1697\ : std_logic;
signal \N__1694\ : std_logic;
signal \N__1691\ : std_logic;
signal \N__1688\ : std_logic;
signal \N__1685\ : std_logic;
signal \N__1682\ : std_logic;
signal \N__1679\ : std_logic;
signal \N__1676\ : std_logic;
signal \N__1673\ : std_logic;
signal \N__1670\ : std_logic;
signal \N__1667\ : std_logic;
signal \N__1664\ : std_logic;
signal \N__1661\ : std_logic;
signal \N__1658\ : std_logic;
signal \N__1655\ : std_logic;
signal \N__1652\ : std_logic;
signal \N__1649\ : std_logic;
signal \N__1646\ : std_logic;
signal \N__1643\ : std_logic;
signal \N__1640\ : std_logic;
signal \N__1637\ : std_logic;
signal \N__1634\ : std_logic;
signal \N__1631\ : std_logic;
signal \N__1628\ : std_logic;
signal \N__1625\ : std_logic;
signal \N__1622\ : std_logic;
signal \N__1619\ : std_logic;
signal \N__1616\ : std_logic;
signal \N__1613\ : std_logic;
signal \N__1610\ : std_logic;
signal \N__1607\ : std_logic;
signal \N__1604\ : std_logic;
signal \N__1601\ : std_logic;
signal \N__1598\ : std_logic;
signal \N__1595\ : std_logic;
signal \N__1592\ : std_logic;
signal \N__1589\ : std_logic;
signal \N__1586\ : std_logic;
signal \N__1583\ : std_logic;
signal \N__1580\ : std_logic;
signal \N__1577\ : std_logic;
signal \N__1574\ : std_logic;
signal \N__1571\ : std_logic;
signal \N__1568\ : std_logic;
signal \N__1565\ : std_logic;
signal \N__1562\ : std_logic;
signal \N__1559\ : std_logic;
signal \N__1556\ : std_logic;
signal \N__1553\ : std_logic;
signal \N__1550\ : std_logic;
signal \N__1547\ : std_logic;
signal \N__1544\ : std_logic;
signal \N__1541\ : std_logic;
signal \N__1538\ : std_logic;
signal \N__1535\ : std_logic;
signal \N__1532\ : std_logic;
signal \N__1529\ : std_logic;
signal \N__1526\ : std_logic;
signal \N__1523\ : std_logic;
signal \N__1520\ : std_logic;
signal \N__1517\ : std_logic;
signal \N__1514\ : std_logic;
signal \N__1511\ : std_logic;
signal \N__1508\ : std_logic;
signal \N__1505\ : std_logic;
signal \N__1502\ : std_logic;
signal \N__1499\ : std_logic;
signal \N__1496\ : std_logic;
signal \N__1493\ : std_logic;
signal \N__1490\ : std_logic;
signal \N__1487\ : std_logic;
signal \N__1484\ : std_logic;
signal \N__1481\ : std_logic;
signal \N__1478\ : std_logic;
signal \N__1475\ : std_logic;
signal \N__1472\ : std_logic;
signal \N__1469\ : std_logic;
signal \N__1466\ : std_logic;
signal \N__1463\ : std_logic;
signal \N__1460\ : std_logic;
signal \N__1457\ : std_logic;
signal \N__1454\ : std_logic;
signal \N__1451\ : std_logic;
signal \N__1448\ : std_logic;
signal \N__1445\ : std_logic;
signal \N__1442\ : std_logic;
signal \N__1439\ : std_logic;
signal \N__1438\ : std_logic;
signal \N__1435\ : std_logic;
signal \N__1432\ : std_logic;
signal \N__1427\ : std_logic;
signal \N__1424\ : std_logic;
signal \N__1421\ : std_logic;
signal \N__1418\ : std_logic;
signal \N__1415\ : std_logic;
signal \N__1412\ : std_logic;
signal \N__1409\ : std_logic;
signal \N__1406\ : std_logic;
signal \N__1403\ : std_logic;
signal \N__1400\ : std_logic;
signal \N__1397\ : std_logic;
signal \N__1394\ : std_logic;
signal \N__1391\ : std_logic;
signal \N__1388\ : std_logic;
signal \N__1385\ : std_logic;
signal \N__1382\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_1\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_2\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_5\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_6\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_3\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_4\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_0\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_10\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_11\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_12\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_13\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_14\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_9\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_7\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_8\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_15\ : std_logic;
signal generated_signal : std_logic;
signal signal_out_c : std_logic;
signal \generator_inst1.REGDYN8_iZ0\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_86\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_87\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_84\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_85\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_9\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_6\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_7\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_8\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_10\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_11\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_12\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_13\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_18\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_14\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_15\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_16\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_17\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_34\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_35\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_36\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_32\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_33\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_37\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_38\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_39\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_40\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_41\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_42\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_43\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_44\ : std_logic;
signal \SELDYN_c\ : std_logic;
signal \SELDYN_c_i\ : std_logic;
signal \RST_N_c\ : std_logic;
signal \RST_N_c_i\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_80\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_81\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_79\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_82\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_83\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_5\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_2\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_3\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_4\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_24\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_23\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_19\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_22\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_20\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_21\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_0\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_1\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_27\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_28\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_29\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_25\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_26\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_30\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_31\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_51\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_52\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_45\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_46\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_47\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_48\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_49\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_50\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_76\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_77\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_78\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_75\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_74\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_73\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_67\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_70\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_68\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_69\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_71\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_72\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_63\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_62\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_60\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_61\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_66\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_64\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_65\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_57\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_58\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_59\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_53\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_54\ : std_logic;
signal \SELSTAT_c\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_55\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_56\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \CLK_c_g\ : std_logic;
signal \SELDYN_c_i_g\ : std_logic;
signal \RST_N_c_i_g\ : std_logic;

signal \CLK_wire\ : std_logic;
signal signal_out_wire : std_logic;
signal \RST_N_wire\ : std_logic;
signal \SELDYN_wire\ : std_logic;
signal \SELSTAT_wire\ : std_logic;

begin
    \CLK_wire\ <= CLK;
    signal_out <= signal_out_wire;
    \RST_N_wire\ <= RST_N;
    \SELDYN_wire\ <= SELDYN;
    \SELSTAT_wire\ <= SELSTAT;

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__2715\,
            GLOBALBUFFEROUTPUT => \CLK_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2717\,
            DIN => \N__2716\,
            DOUT => \N__2715\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2717\,
            PADOUT => \N__2716\,
            PADIN => \N__2715\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \signal_out_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2706\,
            DIN => \N__2705\,
            DOUT => \N__2704\,
            PACKAGEPIN => signal_out_wire
        );

    \signal_out_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2706\,
            PADOUT => \N__2705\,
            PADIN => \N__2704\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1460\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RST_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2697\,
            DIN => \N__2696\,
            DOUT => \N__2695\,
            PACKAGEPIN => \RST_N_wire\
        );

    \RST_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2697\,
            PADOUT => \N__2696\,
            PADIN => \N__2695\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RST_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SELDYN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2688\,
            DIN => \N__2687\,
            DOUT => \N__2686\,
            PACKAGEPIN => \SELDYN_wire\
        );

    \SELDYN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2688\,
            PADOUT => \N__2687\,
            PADIN => \N__2686\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SELDYN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SELSTAT_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2679\,
            DIN => \N__2678\,
            DOUT => \N__2677\,
            PACKAGEPIN => \SELSTAT_wire\
        );

    \SELSTAT_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2679\,
            PADOUT => \N__2678\,
            PADIN => \N__2677\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SELSTAT_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__545\ : InMux
    port map (
            O => \N__2660\,
            I => \N__2657\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__2657\,
            I => \generator_inst1.REGSTATZ0Z_66\
        );

    \I__543\ : InMux
    port map (
            O => \N__2654\,
            I => \N__2651\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__2651\,
            I => \generator_inst1.REGSTATZ0Z_64\
        );

    \I__541\ : InMux
    port map (
            O => \N__2648\,
            I => \N__2645\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__2645\,
            I => \generator_inst1.REGSTATZ0Z_65\
        );

    \I__539\ : InMux
    port map (
            O => \N__2642\,
            I => \N__2639\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__2639\,
            I => \generator_inst1.REGSTATZ0Z_57\
        );

    \I__537\ : InMux
    port map (
            O => \N__2636\,
            I => \N__2633\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__2633\,
            I => \generator_inst1.REGSTATZ0Z_58\
        );

    \I__535\ : InMux
    port map (
            O => \N__2630\,
            I => \N__2627\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__2627\,
            I => \generator_inst1.REGSTATZ0Z_59\
        );

    \I__533\ : InMux
    port map (
            O => \N__2624\,
            I => \N__2621\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__2621\,
            I => \generator_inst1.REGSTATZ0Z_53\
        );

    \I__531\ : InMux
    port map (
            O => \N__2618\,
            I => \N__2615\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__2615\,
            I => \generator_inst1.REGSTATZ0Z_54\
        );

    \I__529\ : InMux
    port map (
            O => \N__2612\,
            I => \N__2560\
        );

    \I__528\ : InMux
    port map (
            O => \N__2611\,
            I => \N__2560\
        );

    \I__527\ : InMux
    port map (
            O => \N__2610\,
            I => \N__2549\
        );

    \I__526\ : InMux
    port map (
            O => \N__2609\,
            I => \N__2549\
        );

    \I__525\ : InMux
    port map (
            O => \N__2608\,
            I => \N__2549\
        );

    \I__524\ : InMux
    port map (
            O => \N__2607\,
            I => \N__2549\
        );

    \I__523\ : InMux
    port map (
            O => \N__2606\,
            I => \N__2549\
        );

    \I__522\ : InMux
    port map (
            O => \N__2605\,
            I => \N__2540\
        );

    \I__521\ : InMux
    port map (
            O => \N__2604\,
            I => \N__2540\
        );

    \I__520\ : InMux
    port map (
            O => \N__2603\,
            I => \N__2540\
        );

    \I__519\ : InMux
    port map (
            O => \N__2602\,
            I => \N__2540\
        );

    \I__518\ : InMux
    port map (
            O => \N__2601\,
            I => \N__2515\
        );

    \I__517\ : InMux
    port map (
            O => \N__2600\,
            I => \N__2515\
        );

    \I__516\ : InMux
    port map (
            O => \N__2599\,
            I => \N__2515\
        );

    \I__515\ : InMux
    port map (
            O => \N__2598\,
            I => \N__2515\
        );

    \I__514\ : InMux
    port map (
            O => \N__2597\,
            I => \N__2515\
        );

    \I__513\ : InMux
    port map (
            O => \N__2596\,
            I => \N__2500\
        );

    \I__512\ : InMux
    port map (
            O => \N__2595\,
            I => \N__2500\
        );

    \I__511\ : InMux
    port map (
            O => \N__2594\,
            I => \N__2500\
        );

    \I__510\ : InMux
    port map (
            O => \N__2593\,
            I => \N__2500\
        );

    \I__509\ : InMux
    port map (
            O => \N__2592\,
            I => \N__2500\
        );

    \I__508\ : InMux
    port map (
            O => \N__2591\,
            I => \N__2500\
        );

    \I__507\ : InMux
    port map (
            O => \N__2590\,
            I => \N__2500\
        );

    \I__506\ : InMux
    port map (
            O => \N__2589\,
            I => \N__2491\
        );

    \I__505\ : InMux
    port map (
            O => \N__2588\,
            I => \N__2491\
        );

    \I__504\ : InMux
    port map (
            O => \N__2587\,
            I => \N__2491\
        );

    \I__503\ : InMux
    port map (
            O => \N__2586\,
            I => \N__2491\
        );

    \I__502\ : InMux
    port map (
            O => \N__2585\,
            I => \N__2476\
        );

    \I__501\ : InMux
    port map (
            O => \N__2584\,
            I => \N__2476\
        );

    \I__500\ : InMux
    port map (
            O => \N__2583\,
            I => \N__2476\
        );

    \I__499\ : InMux
    port map (
            O => \N__2582\,
            I => \N__2476\
        );

    \I__498\ : InMux
    port map (
            O => \N__2581\,
            I => \N__2476\
        );

    \I__497\ : InMux
    port map (
            O => \N__2580\,
            I => \N__2476\
        );

    \I__496\ : InMux
    port map (
            O => \N__2579\,
            I => \N__2476\
        );

    \I__495\ : InMux
    port map (
            O => \N__2578\,
            I => \N__2459\
        );

    \I__494\ : InMux
    port map (
            O => \N__2577\,
            I => \N__2459\
        );

    \I__493\ : InMux
    port map (
            O => \N__2576\,
            I => \N__2459\
        );

    \I__492\ : InMux
    port map (
            O => \N__2575\,
            I => \N__2459\
        );

    \I__491\ : InMux
    port map (
            O => \N__2574\,
            I => \N__2459\
        );

    \I__490\ : InMux
    port map (
            O => \N__2573\,
            I => \N__2459\
        );

    \I__489\ : InMux
    port map (
            O => \N__2572\,
            I => \N__2459\
        );

    \I__488\ : InMux
    port map (
            O => \N__2571\,
            I => \N__2459\
        );

    \I__487\ : InMux
    port map (
            O => \N__2570\,
            I => \N__2446\
        );

    \I__486\ : InMux
    port map (
            O => \N__2569\,
            I => \N__2446\
        );

    \I__485\ : InMux
    port map (
            O => \N__2568\,
            I => \N__2446\
        );

    \I__484\ : InMux
    port map (
            O => \N__2567\,
            I => \N__2446\
        );

    \I__483\ : InMux
    port map (
            O => \N__2566\,
            I => \N__2446\
        );

    \I__482\ : InMux
    port map (
            O => \N__2565\,
            I => \N__2446\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2560\,
            I => \N__2443\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__2549\,
            I => \N__2438\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__2540\,
            I => \N__2438\
        );

    \I__478\ : InMux
    port map (
            O => \N__2539\,
            I => \N__2425\
        );

    \I__477\ : InMux
    port map (
            O => \N__2538\,
            I => \N__2425\
        );

    \I__476\ : InMux
    port map (
            O => \N__2537\,
            I => \N__2425\
        );

    \I__475\ : InMux
    port map (
            O => \N__2536\,
            I => \N__2425\
        );

    \I__474\ : InMux
    port map (
            O => \N__2535\,
            I => \N__2425\
        );

    \I__473\ : InMux
    port map (
            O => \N__2534\,
            I => \N__2425\
        );

    \I__472\ : InMux
    port map (
            O => \N__2533\,
            I => \N__2408\
        );

    \I__471\ : InMux
    port map (
            O => \N__2532\,
            I => \N__2408\
        );

    \I__470\ : InMux
    port map (
            O => \N__2531\,
            I => \N__2408\
        );

    \I__469\ : InMux
    port map (
            O => \N__2530\,
            I => \N__2408\
        );

    \I__468\ : InMux
    port map (
            O => \N__2529\,
            I => \N__2408\
        );

    \I__467\ : InMux
    port map (
            O => \N__2528\,
            I => \N__2408\
        );

    \I__466\ : InMux
    port map (
            O => \N__2527\,
            I => \N__2408\
        );

    \I__465\ : InMux
    port map (
            O => \N__2526\,
            I => \N__2408\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__2515\,
            I => \N__2395\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__2500\,
            I => \N__2395\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__2491\,
            I => \N__2395\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__2476\,
            I => \N__2395\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__2459\,
            I => \N__2395\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__2446\,
            I => \N__2395\
        );

    \I__458\ : Span4Mux_v
    port map (
            O => \N__2443\,
            I => \N__2386\
        );

    \I__457\ : Span4Mux_h
    port map (
            O => \N__2438\,
            I => \N__2386\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__2425\,
            I => \N__2386\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__2408\,
            I => \N__2386\
        );

    \I__454\ : Span4Mux_v
    port map (
            O => \N__2395\,
            I => \N__2361\
        );

    \I__453\ : Span4Mux_v
    port map (
            O => \N__2386\,
            I => \N__2358\
        );

    \I__452\ : InMux
    port map (
            O => \N__2385\,
            I => \N__2345\
        );

    \I__451\ : InMux
    port map (
            O => \N__2384\,
            I => \N__2345\
        );

    \I__450\ : InMux
    port map (
            O => \N__2383\,
            I => \N__2345\
        );

    \I__449\ : InMux
    port map (
            O => \N__2382\,
            I => \N__2345\
        );

    \I__448\ : InMux
    port map (
            O => \N__2381\,
            I => \N__2345\
        );

    \I__447\ : InMux
    port map (
            O => \N__2380\,
            I => \N__2345\
        );

    \I__446\ : InMux
    port map (
            O => \N__2379\,
            I => \N__2328\
        );

    \I__445\ : InMux
    port map (
            O => \N__2378\,
            I => \N__2328\
        );

    \I__444\ : InMux
    port map (
            O => \N__2377\,
            I => \N__2328\
        );

    \I__443\ : InMux
    port map (
            O => \N__2376\,
            I => \N__2328\
        );

    \I__442\ : InMux
    port map (
            O => \N__2375\,
            I => \N__2328\
        );

    \I__441\ : InMux
    port map (
            O => \N__2374\,
            I => \N__2328\
        );

    \I__440\ : InMux
    port map (
            O => \N__2373\,
            I => \N__2328\
        );

    \I__439\ : InMux
    port map (
            O => \N__2372\,
            I => \N__2328\
        );

    \I__438\ : InMux
    port map (
            O => \N__2371\,
            I => \N__2305\
        );

    \I__437\ : InMux
    port map (
            O => \N__2370\,
            I => \N__2305\
        );

    \I__436\ : InMux
    port map (
            O => \N__2369\,
            I => \N__2305\
        );

    \I__435\ : InMux
    port map (
            O => \N__2368\,
            I => \N__2305\
        );

    \I__434\ : InMux
    port map (
            O => \N__2367\,
            I => \N__2305\
        );

    \I__433\ : InMux
    port map (
            O => \N__2366\,
            I => \N__2305\
        );

    \I__432\ : InMux
    port map (
            O => \N__2365\,
            I => \N__2305\
        );

    \I__431\ : InMux
    port map (
            O => \N__2364\,
            I => \N__2305\
        );

    \I__430\ : Sp12to4
    port map (
            O => \N__2361\,
            I => \N__2296\
        );

    \I__429\ : Sp12to4
    port map (
            O => \N__2358\,
            I => \N__2296\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2345\,
            I => \N__2296\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__2328\,
            I => \N__2296\
        );

    \I__426\ : InMux
    port map (
            O => \N__2327\,
            I => \N__2283\
        );

    \I__425\ : InMux
    port map (
            O => \N__2326\,
            I => \N__2283\
        );

    \I__424\ : InMux
    port map (
            O => \N__2325\,
            I => \N__2283\
        );

    \I__423\ : InMux
    port map (
            O => \N__2324\,
            I => \N__2283\
        );

    \I__422\ : InMux
    port map (
            O => \N__2323\,
            I => \N__2283\
        );

    \I__421\ : InMux
    port map (
            O => \N__2322\,
            I => \N__2283\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__2305\,
            I => \SELSTAT_c\
        );

    \I__419\ : Odrv12
    port map (
            O => \N__2296\,
            I => \SELSTAT_c\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__2283\,
            I => \SELSTAT_c\
        );

    \I__417\ : InMux
    port map (
            O => \N__2276\,
            I => \N__2273\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__2273\,
            I => \generator_inst1.REGSTATZ0Z_55\
        );

    \I__415\ : InMux
    port map (
            O => \N__2270\,
            I => \N__2267\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__2267\,
            I => \generator_inst1.REGSTATZ0Z_56\
        );

    \I__413\ : ClkMux
    port map (
            O => \N__2264\,
            I => \N__2213\
        );

    \I__412\ : ClkMux
    port map (
            O => \N__2263\,
            I => \N__2213\
        );

    \I__411\ : ClkMux
    port map (
            O => \N__2262\,
            I => \N__2213\
        );

    \I__410\ : ClkMux
    port map (
            O => \N__2261\,
            I => \N__2213\
        );

    \I__409\ : ClkMux
    port map (
            O => \N__2260\,
            I => \N__2213\
        );

    \I__408\ : ClkMux
    port map (
            O => \N__2259\,
            I => \N__2213\
        );

    \I__407\ : ClkMux
    port map (
            O => \N__2258\,
            I => \N__2213\
        );

    \I__406\ : ClkMux
    port map (
            O => \N__2257\,
            I => \N__2213\
        );

    \I__405\ : ClkMux
    port map (
            O => \N__2256\,
            I => \N__2213\
        );

    \I__404\ : ClkMux
    port map (
            O => \N__2255\,
            I => \N__2213\
        );

    \I__403\ : ClkMux
    port map (
            O => \N__2254\,
            I => \N__2213\
        );

    \I__402\ : ClkMux
    port map (
            O => \N__2253\,
            I => \N__2213\
        );

    \I__401\ : ClkMux
    port map (
            O => \N__2252\,
            I => \N__2213\
        );

    \I__400\ : ClkMux
    port map (
            O => \N__2251\,
            I => \N__2213\
        );

    \I__399\ : ClkMux
    port map (
            O => \N__2250\,
            I => \N__2213\
        );

    \I__398\ : ClkMux
    port map (
            O => \N__2249\,
            I => \N__2213\
        );

    \I__397\ : ClkMux
    port map (
            O => \N__2248\,
            I => \N__2213\
        );

    \I__396\ : GlobalMux
    port map (
            O => \N__2213\,
            I => \N__2210\
        );

    \I__395\ : gio2CtrlBuf
    port map (
            O => \N__2210\,
            I => \CLK_c_g\
        );

    \I__394\ : CEMux
    port map (
            O => \N__2207\,
            I => \N__2165\
        );

    \I__393\ : CEMux
    port map (
            O => \N__2206\,
            I => \N__2165\
        );

    \I__392\ : CEMux
    port map (
            O => \N__2205\,
            I => \N__2165\
        );

    \I__391\ : CEMux
    port map (
            O => \N__2204\,
            I => \N__2165\
        );

    \I__390\ : CEMux
    port map (
            O => \N__2203\,
            I => \N__2165\
        );

    \I__389\ : CEMux
    port map (
            O => \N__2202\,
            I => \N__2165\
        );

    \I__388\ : CEMux
    port map (
            O => \N__2201\,
            I => \N__2165\
        );

    \I__387\ : CEMux
    port map (
            O => \N__2200\,
            I => \N__2165\
        );

    \I__386\ : CEMux
    port map (
            O => \N__2199\,
            I => \N__2165\
        );

    \I__385\ : CEMux
    port map (
            O => \N__2198\,
            I => \N__2165\
        );

    \I__384\ : CEMux
    port map (
            O => \N__2197\,
            I => \N__2165\
        );

    \I__383\ : CEMux
    port map (
            O => \N__2196\,
            I => \N__2165\
        );

    \I__382\ : CEMux
    port map (
            O => \N__2195\,
            I => \N__2165\
        );

    \I__381\ : CEMux
    port map (
            O => \N__2194\,
            I => \N__2165\
        );

    \I__380\ : GlobalMux
    port map (
            O => \N__2165\,
            I => \N__2162\
        );

    \I__379\ : gio2CtrlBuf
    port map (
            O => \N__2162\,
            I => \SELDYN_c_i_g\
        );

    \I__378\ : SRMux
    port map (
            O => \N__2159\,
            I => \N__2108\
        );

    \I__377\ : SRMux
    port map (
            O => \N__2158\,
            I => \N__2108\
        );

    \I__376\ : SRMux
    port map (
            O => \N__2157\,
            I => \N__2108\
        );

    \I__375\ : SRMux
    port map (
            O => \N__2156\,
            I => \N__2108\
        );

    \I__374\ : SRMux
    port map (
            O => \N__2155\,
            I => \N__2108\
        );

    \I__373\ : SRMux
    port map (
            O => \N__2154\,
            I => \N__2108\
        );

    \I__372\ : SRMux
    port map (
            O => \N__2153\,
            I => \N__2108\
        );

    \I__371\ : SRMux
    port map (
            O => \N__2152\,
            I => \N__2108\
        );

    \I__370\ : SRMux
    port map (
            O => \N__2151\,
            I => \N__2108\
        );

    \I__369\ : SRMux
    port map (
            O => \N__2150\,
            I => \N__2108\
        );

    \I__368\ : SRMux
    port map (
            O => \N__2149\,
            I => \N__2108\
        );

    \I__367\ : SRMux
    port map (
            O => \N__2148\,
            I => \N__2108\
        );

    \I__366\ : SRMux
    port map (
            O => \N__2147\,
            I => \N__2108\
        );

    \I__365\ : SRMux
    port map (
            O => \N__2146\,
            I => \N__2108\
        );

    \I__364\ : SRMux
    port map (
            O => \N__2145\,
            I => \N__2108\
        );

    \I__363\ : SRMux
    port map (
            O => \N__2144\,
            I => \N__2108\
        );

    \I__362\ : SRMux
    port map (
            O => \N__2143\,
            I => \N__2108\
        );

    \I__361\ : GlobalMux
    port map (
            O => \N__2108\,
            I => \N__2105\
        );

    \I__360\ : gio2CtrlBuf
    port map (
            O => \N__2105\,
            I => \RST_N_c_i_g\
        );

    \I__359\ : InMux
    port map (
            O => \N__2102\,
            I => \N__2099\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2099\,
            I => \generator_inst1.REGSTATZ0Z_67\
        );

    \I__357\ : InMux
    port map (
            O => \N__2096\,
            I => \N__2093\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2093\,
            I => \generator_inst1.REGSTATZ0Z_70\
        );

    \I__355\ : InMux
    port map (
            O => \N__2090\,
            I => \N__2087\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__2087\,
            I => \generator_inst1.REGSTATZ0Z_68\
        );

    \I__353\ : InMux
    port map (
            O => \N__2084\,
            I => \N__2081\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__2081\,
            I => \generator_inst1.REGSTATZ0Z_69\
        );

    \I__351\ : InMux
    port map (
            O => \N__2078\,
            I => \N__2075\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2075\,
            I => \generator_inst1.REGSTATZ0Z_71\
        );

    \I__349\ : InMux
    port map (
            O => \N__2072\,
            I => \N__2069\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__2069\,
            I => \generator_inst1.REGSTATZ0Z_72\
        );

    \I__347\ : InMux
    port map (
            O => \N__2066\,
            I => \N__2063\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2063\,
            I => \generator_inst1.REGSTATZ0Z_63\
        );

    \I__345\ : InMux
    port map (
            O => \N__2060\,
            I => \N__2057\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__2057\,
            I => \generator_inst1.REGSTATZ0Z_62\
        );

    \I__343\ : InMux
    port map (
            O => \N__2054\,
            I => \N__2051\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2051\,
            I => \generator_inst1.REGSTATZ0Z_60\
        );

    \I__341\ : InMux
    port map (
            O => \N__2048\,
            I => \N__2045\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2045\,
            I => \generator_inst1.REGSTATZ0Z_61\
        );

    \I__339\ : InMux
    port map (
            O => \N__2042\,
            I => \N__2039\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2039\,
            I => \generator_inst1.REGSTATZ0Z_49\
        );

    \I__337\ : InMux
    port map (
            O => \N__2036\,
            I => \N__2033\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2033\,
            I => \generator_inst1.REGSTATZ0Z_50\
        );

    \I__335\ : InMux
    port map (
            O => \N__2030\,
            I => \N__2027\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2027\,
            I => \generator_inst1.REGSTATZ0Z_76\
        );

    \I__333\ : InMux
    port map (
            O => \N__2024\,
            I => \N__2021\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2021\,
            I => \generator_inst1.REGSTATZ0Z_77\
        );

    \I__331\ : InMux
    port map (
            O => \N__2018\,
            I => \N__2015\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2015\,
            I => \generator_inst1.REGSTATZ0Z_78\
        );

    \I__329\ : InMux
    port map (
            O => \N__2012\,
            I => \N__2009\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2009\,
            I => \generator_inst1.REGSTATZ0Z_75\
        );

    \I__327\ : InMux
    port map (
            O => \N__2006\,
            I => \N__2003\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__2003\,
            I => \generator_inst1.REGSTATZ0Z_74\
        );

    \I__325\ : InMux
    port map (
            O => \N__2000\,
            I => \N__1997\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__1997\,
            I => \generator_inst1.REGSTATZ0Z_73\
        );

    \I__323\ : InMux
    port map (
            O => \N__1994\,
            I => \N__1991\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__1991\,
            I => \generator_inst1.REGSTATZ0Z_25\
        );

    \I__321\ : InMux
    port map (
            O => \N__1988\,
            I => \N__1985\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__1985\,
            I => \generator_inst1.REGSTATZ0Z_26\
        );

    \I__319\ : InMux
    port map (
            O => \N__1982\,
            I => \N__1979\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__1979\,
            I => \generator_inst1.REGSTATZ0Z_30\
        );

    \I__317\ : InMux
    port map (
            O => \N__1976\,
            I => \N__1973\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__1973\,
            I => \generator_inst1.REGSTATZ0Z_31\
        );

    \I__315\ : InMux
    port map (
            O => \N__1970\,
            I => \N__1967\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__1967\,
            I => \generator_inst1.REGSTATZ0Z_51\
        );

    \I__313\ : InMux
    port map (
            O => \N__1964\,
            I => \N__1961\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__1961\,
            I => \generator_inst1.REGSTATZ0Z_52\
        );

    \I__311\ : InMux
    port map (
            O => \N__1958\,
            I => \N__1955\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__1955\,
            I => \generator_inst1.REGSTATZ0Z_45\
        );

    \I__309\ : InMux
    port map (
            O => \N__1952\,
            I => \N__1949\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__1949\,
            I => \generator_inst1.REGSTATZ0Z_46\
        );

    \I__307\ : InMux
    port map (
            O => \N__1946\,
            I => \N__1943\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__1943\,
            I => \generator_inst1.REGSTATZ0Z_47\
        );

    \I__305\ : InMux
    port map (
            O => \N__1940\,
            I => \N__1937\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__1937\,
            I => \generator_inst1.REGSTATZ0Z_48\
        );

    \I__303\ : InMux
    port map (
            O => \N__1934\,
            I => \N__1931\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__1931\,
            I => \generator_inst1.REGSTATZ0Z_19\
        );

    \I__301\ : InMux
    port map (
            O => \N__1928\,
            I => \N__1925\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__1925\,
            I => \generator_inst1.REGSTATZ0Z_22\
        );

    \I__299\ : InMux
    port map (
            O => \N__1922\,
            I => \N__1919\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__1919\,
            I => \generator_inst1.REGSTATZ0Z_20\
        );

    \I__297\ : InMux
    port map (
            O => \N__1916\,
            I => \N__1913\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__1913\,
            I => \generator_inst1.REGSTATZ0Z_21\
        );

    \I__295\ : InMux
    port map (
            O => \N__1910\,
            I => \N__1907\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__1907\,
            I => \generator_inst1.REGSTATZ0Z_0\
        );

    \I__293\ : InMux
    port map (
            O => \N__1904\,
            I => \N__1901\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__1901\,
            I => \generator_inst1.REGSTATZ0Z_1\
        );

    \I__291\ : InMux
    port map (
            O => \N__1898\,
            I => \N__1895\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__1895\,
            I => \generator_inst1.REGSTATZ0Z_27\
        );

    \I__289\ : InMux
    port map (
            O => \N__1892\,
            I => \N__1889\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__1889\,
            I => \generator_inst1.REGSTATZ0Z_28\
        );

    \I__287\ : InMux
    port map (
            O => \N__1886\,
            I => \N__1883\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__1883\,
            I => \generator_inst1.REGSTATZ0Z_29\
        );

    \I__285\ : InMux
    port map (
            O => \N__1880\,
            I => \N__1877\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__1877\,
            I => \generator_inst1.REGSTATZ0Z_79\
        );

    \I__283\ : InMux
    port map (
            O => \N__1874\,
            I => \N__1871\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__1871\,
            I => \generator_inst1.REGSTATZ0Z_82\
        );

    \I__281\ : InMux
    port map (
            O => \N__1868\,
            I => \N__1865\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__1865\,
            I => \generator_inst1.REGSTATZ0Z_83\
        );

    \I__279\ : InMux
    port map (
            O => \N__1862\,
            I => \N__1859\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__1859\,
            I => \generator_inst1.REGSTATZ0Z_5\
        );

    \I__277\ : InMux
    port map (
            O => \N__1856\,
            I => \N__1853\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__1853\,
            I => \generator_inst1.REGSTATZ0Z_2\
        );

    \I__275\ : InMux
    port map (
            O => \N__1850\,
            I => \N__1847\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__1847\,
            I => \generator_inst1.REGSTATZ0Z_3\
        );

    \I__273\ : InMux
    port map (
            O => \N__1844\,
            I => \N__1841\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__1841\,
            I => \generator_inst1.REGSTATZ0Z_4\
        );

    \I__271\ : InMux
    port map (
            O => \N__1838\,
            I => \N__1835\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__1835\,
            I => \generator_inst1.REGSTATZ0Z_24\
        );

    \I__269\ : InMux
    port map (
            O => \N__1832\,
            I => \N__1829\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__1829\,
            I => \generator_inst1.REGSTATZ0Z_23\
        );

    \I__267\ : InMux
    port map (
            O => \N__1826\,
            I => \N__1823\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__1823\,
            I => \generator_inst1.REGSTATZ0Z_40\
        );

    \I__265\ : InMux
    port map (
            O => \N__1820\,
            I => \N__1817\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__1817\,
            I => \generator_inst1.REGSTATZ0Z_41\
        );

    \I__263\ : InMux
    port map (
            O => \N__1814\,
            I => \N__1811\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__1811\,
            I => \generator_inst1.REGSTATZ0Z_42\
        );

    \I__261\ : InMux
    port map (
            O => \N__1808\,
            I => \N__1805\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__1805\,
            I => \generator_inst1.REGSTATZ0Z_43\
        );

    \I__259\ : InMux
    port map (
            O => \N__1802\,
            I => \N__1799\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__1799\,
            I => \generator_inst1.REGSTATZ0Z_44\
        );

    \I__257\ : InMux
    port map (
            O => \N__1796\,
            I => \N__1793\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__1793\,
            I => \N__1790\
        );

    \I__255\ : Span4Mux_v
    port map (
            O => \N__1790\,
            I => \N__1769\
        );

    \I__254\ : InMux
    port map (
            O => \N__1789\,
            I => \N__1764\
        );

    \I__253\ : InMux
    port map (
            O => \N__1788\,
            I => \N__1764\
        );

    \I__252\ : InMux
    port map (
            O => \N__1787\,
            I => \N__1747\
        );

    \I__251\ : InMux
    port map (
            O => \N__1786\,
            I => \N__1747\
        );

    \I__250\ : InMux
    port map (
            O => \N__1785\,
            I => \N__1747\
        );

    \I__249\ : InMux
    port map (
            O => \N__1784\,
            I => \N__1747\
        );

    \I__248\ : InMux
    port map (
            O => \N__1783\,
            I => \N__1747\
        );

    \I__247\ : InMux
    port map (
            O => \N__1782\,
            I => \N__1747\
        );

    \I__246\ : InMux
    port map (
            O => \N__1781\,
            I => \N__1747\
        );

    \I__245\ : InMux
    port map (
            O => \N__1780\,
            I => \N__1747\
        );

    \I__244\ : InMux
    port map (
            O => \N__1779\,
            I => \N__1730\
        );

    \I__243\ : InMux
    port map (
            O => \N__1778\,
            I => \N__1730\
        );

    \I__242\ : InMux
    port map (
            O => \N__1777\,
            I => \N__1730\
        );

    \I__241\ : InMux
    port map (
            O => \N__1776\,
            I => \N__1730\
        );

    \I__240\ : InMux
    port map (
            O => \N__1775\,
            I => \N__1730\
        );

    \I__239\ : InMux
    port map (
            O => \N__1774\,
            I => \N__1730\
        );

    \I__238\ : InMux
    port map (
            O => \N__1773\,
            I => \N__1730\
        );

    \I__237\ : InMux
    port map (
            O => \N__1772\,
            I => \N__1730\
        );

    \I__236\ : Span4Mux_v
    port map (
            O => \N__1769\,
            I => \N__1721\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__1764\,
            I => \N__1721\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__1747\,
            I => \N__1721\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__1730\,
            I => \N__1721\
        );

    \I__232\ : Span4Mux_v
    port map (
            O => \N__1721\,
            I => \N__1718\
        );

    \I__231\ : Span4Mux_v
    port map (
            O => \N__1718\,
            I => \N__1715\
        );

    \I__230\ : Odrv4
    port map (
            O => \N__1715\,
            I => \SELDYN_c\
        );

    \I__229\ : IoInMux
    port map (
            O => \N__1712\,
            I => \N__1709\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__1709\,
            I => \SELDYN_c_i\
        );

    \I__227\ : InMux
    port map (
            O => \N__1706\,
            I => \N__1703\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__1703\,
            I => \N__1700\
        );

    \I__225\ : Span4Mux_v
    port map (
            O => \N__1700\,
            I => \N__1697\
        );

    \I__224\ : Span4Mux_v
    port map (
            O => \N__1697\,
            I => \N__1694\
        );

    \I__223\ : Odrv4
    port map (
            O => \N__1694\,
            I => \RST_N_c\
        );

    \I__222\ : IoInMux
    port map (
            O => \N__1691\,
            I => \N__1688\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__1688\,
            I => \N__1685\
        );

    \I__220\ : IoSpan4Mux
    port map (
            O => \N__1685\,
            I => \N__1682\
        );

    \I__219\ : Odrv4
    port map (
            O => \N__1682\,
            I => \RST_N_c_i\
        );

    \I__218\ : InMux
    port map (
            O => \N__1679\,
            I => \N__1676\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__1676\,
            I => \generator_inst1.REGSTATZ0Z_80\
        );

    \I__216\ : InMux
    port map (
            O => \N__1673\,
            I => \N__1670\
        );

    \I__215\ : LocalMux
    port map (
            O => \N__1670\,
            I => \generator_inst1.REGSTATZ0Z_81\
        );

    \I__214\ : InMux
    port map (
            O => \N__1667\,
            I => \N__1664\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__1664\,
            I => \generator_inst1.REGSTATZ0Z_34\
        );

    \I__212\ : InMux
    port map (
            O => \N__1661\,
            I => \N__1658\
        );

    \I__211\ : LocalMux
    port map (
            O => \N__1658\,
            I => \generator_inst1.REGSTATZ0Z_35\
        );

    \I__210\ : InMux
    port map (
            O => \N__1655\,
            I => \N__1652\
        );

    \I__209\ : LocalMux
    port map (
            O => \N__1652\,
            I => \generator_inst1.REGSTATZ0Z_36\
        );

    \I__208\ : InMux
    port map (
            O => \N__1649\,
            I => \N__1646\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__1646\,
            I => \generator_inst1.REGSTATZ0Z_32\
        );

    \I__206\ : InMux
    port map (
            O => \N__1643\,
            I => \N__1640\
        );

    \I__205\ : LocalMux
    port map (
            O => \N__1640\,
            I => \generator_inst1.REGSTATZ0Z_33\
        );

    \I__204\ : InMux
    port map (
            O => \N__1637\,
            I => \N__1634\
        );

    \I__203\ : LocalMux
    port map (
            O => \N__1634\,
            I => \generator_inst1.REGSTATZ0Z_37\
        );

    \I__202\ : InMux
    port map (
            O => \N__1631\,
            I => \N__1628\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__1628\,
            I => \generator_inst1.REGSTATZ0Z_38\
        );

    \I__200\ : InMux
    port map (
            O => \N__1625\,
            I => \N__1622\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__1622\,
            I => \generator_inst1.REGSTATZ0Z_39\
        );

    \I__198\ : InMux
    port map (
            O => \N__1619\,
            I => \N__1616\
        );

    \I__197\ : LocalMux
    port map (
            O => \N__1616\,
            I => \generator_inst1.REGSTATZ0Z_10\
        );

    \I__196\ : InMux
    port map (
            O => \N__1613\,
            I => \N__1610\
        );

    \I__195\ : LocalMux
    port map (
            O => \N__1610\,
            I => \generator_inst1.REGSTATZ0Z_11\
        );

    \I__194\ : InMux
    port map (
            O => \N__1607\,
            I => \N__1604\
        );

    \I__193\ : LocalMux
    port map (
            O => \N__1604\,
            I => \generator_inst1.REGSTATZ0Z_12\
        );

    \I__192\ : InMux
    port map (
            O => \N__1601\,
            I => \N__1598\
        );

    \I__191\ : LocalMux
    port map (
            O => \N__1598\,
            I => \generator_inst1.REGSTATZ0Z_13\
        );

    \I__190\ : InMux
    port map (
            O => \N__1595\,
            I => \N__1592\
        );

    \I__189\ : LocalMux
    port map (
            O => \N__1592\,
            I => \generator_inst1.REGSTATZ0Z_18\
        );

    \I__188\ : InMux
    port map (
            O => \N__1589\,
            I => \N__1586\
        );

    \I__187\ : LocalMux
    port map (
            O => \N__1586\,
            I => \generator_inst1.REGSTATZ0Z_14\
        );

    \I__186\ : InMux
    port map (
            O => \N__1583\,
            I => \N__1580\
        );

    \I__185\ : LocalMux
    port map (
            O => \N__1580\,
            I => \generator_inst1.REGSTATZ0Z_15\
        );

    \I__184\ : InMux
    port map (
            O => \N__1577\,
            I => \N__1574\
        );

    \I__183\ : LocalMux
    port map (
            O => \N__1574\,
            I => \generator_inst1.REGSTATZ0Z_16\
        );

    \I__182\ : InMux
    port map (
            O => \N__1571\,
            I => \N__1568\
        );

    \I__181\ : LocalMux
    port map (
            O => \N__1568\,
            I => \generator_inst1.REGSTATZ0Z_17\
        );

    \I__180\ : InMux
    port map (
            O => \N__1565\,
            I => \N__1562\
        );

    \I__179\ : LocalMux
    port map (
            O => \N__1562\,
            I => \generator_inst1.REGSTATZ0Z_86\
        );

    \I__178\ : CascadeMux
    port map (
            O => \N__1559\,
            I => \N__1556\
        );

    \I__177\ : InMux
    port map (
            O => \N__1556\,
            I => \N__1553\
        );

    \I__176\ : LocalMux
    port map (
            O => \N__1553\,
            I => \generator_inst1.REGSTATZ0Z_87\
        );

    \I__175\ : InMux
    port map (
            O => \N__1550\,
            I => \N__1547\
        );

    \I__174\ : LocalMux
    port map (
            O => \N__1547\,
            I => \generator_inst1.REGSTATZ0Z_84\
        );

    \I__173\ : InMux
    port map (
            O => \N__1544\,
            I => \N__1541\
        );

    \I__172\ : LocalMux
    port map (
            O => \N__1541\,
            I => \generator_inst1.REGSTATZ0Z_85\
        );

    \I__171\ : InMux
    port map (
            O => \N__1538\,
            I => \N__1535\
        );

    \I__170\ : LocalMux
    port map (
            O => \N__1535\,
            I => \generator_inst1.REGSTATZ0Z_9\
        );

    \I__169\ : InMux
    port map (
            O => \N__1532\,
            I => \N__1529\
        );

    \I__168\ : LocalMux
    port map (
            O => \N__1529\,
            I => \generator_inst1.REGSTATZ0Z_6\
        );

    \I__167\ : InMux
    port map (
            O => \N__1526\,
            I => \N__1523\
        );

    \I__166\ : LocalMux
    port map (
            O => \N__1523\,
            I => \generator_inst1.REGSTATZ0Z_7\
        );

    \I__165\ : InMux
    port map (
            O => \N__1520\,
            I => \N__1517\
        );

    \I__164\ : LocalMux
    port map (
            O => \N__1517\,
            I => \generator_inst1.REGSTATZ0Z_8\
        );

    \I__163\ : InMux
    port map (
            O => \N__1514\,
            I => \N__1511\
        );

    \I__162\ : LocalMux
    port map (
            O => \N__1511\,
            I => \generator_inst1.REGDYNZ0Z_11\
        );

    \I__161\ : InMux
    port map (
            O => \N__1508\,
            I => \N__1505\
        );

    \I__160\ : LocalMux
    port map (
            O => \N__1505\,
            I => \generator_inst1.REGDYNZ0Z_12\
        );

    \I__159\ : InMux
    port map (
            O => \N__1502\,
            I => \N__1499\
        );

    \I__158\ : LocalMux
    port map (
            O => \N__1499\,
            I => \generator_inst1.REGDYNZ0Z_13\
        );

    \I__157\ : InMux
    port map (
            O => \N__1496\,
            I => \N__1493\
        );

    \I__156\ : LocalMux
    port map (
            O => \N__1493\,
            I => \generator_inst1.REGDYNZ0Z_14\
        );

    \I__155\ : InMux
    port map (
            O => \N__1490\,
            I => \N__1487\
        );

    \I__154\ : LocalMux
    port map (
            O => \N__1487\,
            I => \generator_inst1.REGDYNZ0Z_9\
        );

    \I__153\ : InMux
    port map (
            O => \N__1484\,
            I => \N__1481\
        );

    \I__152\ : LocalMux
    port map (
            O => \N__1481\,
            I => \generator_inst1.REGDYNZ0Z_7\
        );

    \I__151\ : InMux
    port map (
            O => \N__1478\,
            I => \N__1475\
        );

    \I__150\ : LocalMux
    port map (
            O => \N__1475\,
            I => \generator_inst1.REGDYNZ0Z_8\
        );

    \I__149\ : InMux
    port map (
            O => \N__1472\,
            I => \N__1469\
        );

    \I__148\ : LocalMux
    port map (
            O => \N__1469\,
            I => \generator_inst1.REGDYNZ0Z_15\
        );

    \I__147\ : InMux
    port map (
            O => \N__1466\,
            I => \N__1463\
        );

    \I__146\ : LocalMux
    port map (
            O => \N__1463\,
            I => generated_signal
        );

    \I__145\ : IoInMux
    port map (
            O => \N__1460\,
            I => \N__1457\
        );

    \I__144\ : LocalMux
    port map (
            O => \N__1457\,
            I => \N__1454\
        );

    \I__143\ : Span4Mux_s1_h
    port map (
            O => \N__1454\,
            I => \N__1451\
        );

    \I__142\ : Span4Mux_v
    port map (
            O => \N__1451\,
            I => \N__1448\
        );

    \I__141\ : Odrv4
    port map (
            O => \N__1448\,
            I => signal_out_c
        );

    \I__140\ : CEMux
    port map (
            O => \N__1445\,
            I => \N__1442\
        );

    \I__139\ : LocalMux
    port map (
            O => \N__1442\,
            I => \N__1439\
        );

    \I__138\ : Sp12to4
    port map (
            O => \N__1439\,
            I => \N__1435\
        );

    \I__137\ : CEMux
    port map (
            O => \N__1438\,
            I => \N__1432\
        );

    \I__136\ : Odrv12
    port map (
            O => \N__1435\,
            I => \generator_inst1.REGDYN8_iZ0\
        );

    \I__135\ : LocalMux
    port map (
            O => \N__1432\,
            I => \generator_inst1.REGDYN8_iZ0\
        );

    \I__134\ : InMux
    port map (
            O => \N__1427\,
            I => \N__1424\
        );

    \I__133\ : LocalMux
    port map (
            O => \N__1424\,
            I => \generator_inst1.REGDYNZ0Z_1\
        );

    \I__132\ : InMux
    port map (
            O => \N__1421\,
            I => \N__1418\
        );

    \I__131\ : LocalMux
    port map (
            O => \N__1418\,
            I => \generator_inst1.REGDYNZ0Z_2\
        );

    \I__130\ : InMux
    port map (
            O => \N__1415\,
            I => \N__1412\
        );

    \I__129\ : LocalMux
    port map (
            O => \N__1412\,
            I => \generator_inst1.REGDYNZ0Z_5\
        );

    \I__128\ : InMux
    port map (
            O => \N__1409\,
            I => \N__1406\
        );

    \I__127\ : LocalMux
    port map (
            O => \N__1406\,
            I => \generator_inst1.REGDYNZ0Z_6\
        );

    \I__126\ : InMux
    port map (
            O => \N__1403\,
            I => \N__1400\
        );

    \I__125\ : LocalMux
    port map (
            O => \N__1400\,
            I => \generator_inst1.REGDYNZ0Z_3\
        );

    \I__124\ : InMux
    port map (
            O => \N__1397\,
            I => \N__1394\
        );

    \I__123\ : LocalMux
    port map (
            O => \N__1394\,
            I => \generator_inst1.REGDYNZ0Z_4\
        );

    \I__122\ : InMux
    port map (
            O => \N__1391\,
            I => \N__1388\
        );

    \I__121\ : LocalMux
    port map (
            O => \N__1388\,
            I => \generator_inst1.REGDYNZ0Z_0\
        );

    \I__120\ : InMux
    port map (
            O => \N__1385\,
            I => \N__1382\
        );

    \I__119\ : LocalMux
    port map (
            O => \N__1382\,
            I => \generator_inst1.REGDYNZ0Z_10\
        );

    \RST_N_ibuf_RNIBJGC_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__1691\,
            GLOBALBUFFEROUTPUT => \RST_N_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \SELDYN_ibuf_RNIKHL3_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__1712\,
            GLOBALBUFFEROUTPUT => \SELDYN_c_i_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \generator_inst1.REGDYN_2_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__1774\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1427\,
            lcout => \generator_inst1.REGDYNZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2264\,
            ce => \N__1445\,
            sr => \N__2159\
        );

    \generator_inst1.REGDYN_1_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1773\,
            in2 => \_gnd_net_\,
            in3 => \N__1391\,
            lcout => \generator_inst1.REGDYNZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2264\,
            ce => \N__1445\,
            sr => \N__2159\
        );

    \generator_inst1.REGDYN_3_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__1775\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1421\,
            lcout => \generator_inst1.REGDYNZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2264\,
            ce => \N__1445\,
            sr => \N__2159\
        );

    \generator_inst1.REGDYN_7_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1779\,
            in2 => \_gnd_net_\,
            in3 => \N__1409\,
            lcout => \generator_inst1.REGDYNZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2264\,
            ce => \N__1445\,
            sr => \N__2159\
        );

    \generator_inst1.REGDYN_5_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__1777\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1397\,
            lcout => \generator_inst1.REGDYNZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2264\,
            ce => \N__1445\,
            sr => \N__2159\
        );

    \generator_inst1.REGDYN_6_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1778\,
            in2 => \_gnd_net_\,
            in3 => \N__1415\,
            lcout => \generator_inst1.REGDYNZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2264\,
            ce => \N__1445\,
            sr => \N__2159\
        );

    \generator_inst1.REGDYN_4_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__1776\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1403\,
            lcout => \generator_inst1.REGDYNZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2264\,
            ce => \N__1445\,
            sr => \N__2159\
        );

    \generator_inst1.REGDYN_0_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1772\,
            lcout => \generator_inst1.REGDYNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2264\,
            ce => \N__1445\,
            sr => \N__2159\
        );

    \generator_inst1.REGDYN_11_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1781\,
            in2 => \_gnd_net_\,
            in3 => \N__1385\,
            lcout => \generator_inst1.REGDYNZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2263\,
            ce => \N__1438\,
            sr => \N__2158\
        );

    \generator_inst1.REGDYN_10_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__1780\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1490\,
            lcout => \generator_inst1.REGDYNZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2263\,
            ce => \N__1438\,
            sr => \N__2158\
        );

    \generator_inst1.REGDYN_12_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1782\,
            in2 => \_gnd_net_\,
            in3 => \N__1514\,
            lcout => \generator_inst1.REGDYNZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2263\,
            ce => \N__1438\,
            sr => \N__2158\
        );

    \generator_inst1.REGDYN_13_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__1783\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1508\,
            lcout => \generator_inst1.REGDYNZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2263\,
            ce => \N__1438\,
            sr => \N__2158\
        );

    \generator_inst1.REGDYN_14_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1784\,
            in2 => \_gnd_net_\,
            in3 => \N__1502\,
            lcout => \generator_inst1.REGDYNZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2263\,
            ce => \N__1438\,
            sr => \N__2158\
        );

    \generator_inst1.REGDYN_15_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__1785\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1496\,
            lcout => \generator_inst1.REGDYNZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2263\,
            ce => \N__1438\,
            sr => \N__2158\
        );

    \generator_inst1.REGDYN_9_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1787\,
            in2 => \_gnd_net_\,
            in3 => \N__1478\,
            lcout => \generator_inst1.REGDYNZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2263\,
            ce => \N__1438\,
            sr => \N__2158\
        );

    \generator_inst1.REGDYN_8_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__1786\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1484\,
            lcout => \generator_inst1.REGDYNZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2263\,
            ce => \N__1438\,
            sr => \N__2158\
        );

    \generator_inst1.signal_out_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110001001000000"
        )
    port map (
            in0 => \N__2612\,
            in1 => \N__1789\,
            in2 => \N__1559\,
            in3 => \N__1472\,
            lcout => generated_signal,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2260\,
            ce => 'H',
            sr => \N__2155\
        );

    \receptor_inst1.signal_out_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1466\,
            lcout => signal_out_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2260\,
            ce => 'H',
            sr => \N__2155\
        );

    \generator_inst1.REGDYN8_i_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__2611\,
            in1 => \N__1788\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \generator_inst1.REGDYN8_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.REGSTAT_86_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2604\,
            in2 => \_gnd_net_\,
            in3 => \N__1544\,
            lcout => \generator_inst1.REGSTATZ0Z_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2257\,
            ce => \N__2203\,
            sr => \N__2152\
        );

    \generator_inst1.REGSTAT_87_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2605\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1565\,
            lcout => \generator_inst1.REGSTATZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2257\,
            ce => \N__2203\,
            sr => \N__2152\
        );

    \generator_inst1.REGSTAT_84_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2602\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1868\,
            lcout => \generator_inst1.REGSTATZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2257\,
            ce => \N__2203\,
            sr => \N__2152\
        );

    \generator_inst1.REGSTAT_85_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2603\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1550\,
            lcout => \generator_inst1.REGSTATZ0Z_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2257\,
            ce => \N__2203\,
            sr => \N__2152\
        );

    \generator_inst1.REGSTAT_10_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2534\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1538\,
            lcout => \generator_inst1.REGSTATZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2254\,
            ce => \N__2200\,
            sr => \N__2149\
        );

    \generator_inst1.REGSTAT_7_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2537\,
            in2 => \_gnd_net_\,
            in3 => \N__1532\,
            lcout => \generator_inst1.REGSTATZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2254\,
            ce => \N__2200\,
            sr => \N__2149\
        );

    \generator_inst1.REGSTAT_9_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2539\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1520\,
            lcout => \generator_inst1.REGSTATZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2254\,
            ce => \N__2200\,
            sr => \N__2149\
        );

    \generator_inst1.REGSTAT_6_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2536\,
            in2 => \_gnd_net_\,
            in3 => \N__1862\,
            lcout => \generator_inst1.REGSTATZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2254\,
            ce => \N__2200\,
            sr => \N__2149\
        );

    \generator_inst1.REGSTAT_8_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2538\,
            in2 => \_gnd_net_\,
            in3 => \N__1526\,
            lcout => \generator_inst1.REGSTATZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2254\,
            ce => \N__2200\,
            sr => \N__2149\
        );

    \generator_inst1.REGSTAT_11_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2535\,
            in2 => \_gnd_net_\,
            in3 => \N__1619\,
            lcout => \generator_inst1.REGSTATZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2254\,
            ce => \N__2200\,
            sr => \N__2149\
        );

    \generator_inst1.REGSTAT_19_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2533\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1595\,
            lcout => \generator_inst1.REGSTATZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2251\,
            ce => \N__2197\,
            sr => \N__2147\
        );

    \generator_inst1.REGSTAT_12_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2526\,
            in2 => \_gnd_net_\,
            in3 => \N__1613\,
            lcout => \generator_inst1.REGSTATZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2251\,
            ce => \N__2197\,
            sr => \N__2147\
        );

    \generator_inst1.REGSTAT_14_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1601\,
            lcout => \generator_inst1.REGSTATZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2251\,
            ce => \N__2197\,
            sr => \N__2147\
        );

    \generator_inst1.REGSTAT_13_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2527\,
            in2 => \_gnd_net_\,
            in3 => \N__1607\,
            lcout => \generator_inst1.REGSTATZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2251\,
            ce => \N__2197\,
            sr => \N__2147\
        );

    \generator_inst1.REGSTAT_18_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2532\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1571\,
            lcout => \generator_inst1.REGSTATZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2251\,
            ce => \N__2197\,
            sr => \N__2147\
        );

    \generator_inst1.REGSTAT_15_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2529\,
            in2 => \_gnd_net_\,
            in3 => \N__1589\,
            lcout => \generator_inst1.REGSTATZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2251\,
            ce => \N__2197\,
            sr => \N__2147\
        );

    \generator_inst1.REGSTAT_16_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2530\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1583\,
            lcout => \generator_inst1.REGSTATZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2251\,
            ce => \N__2197\,
            sr => \N__2147\
        );

    \generator_inst1.REGSTAT_17_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2531\,
            in2 => \_gnd_net_\,
            in3 => \N__1577\,
            lcout => \generator_inst1.REGSTATZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2251\,
            ce => \N__2197\,
            sr => \N__2147\
        );

    \generator_inst1.REGSTAT_32_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2364\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1976\,
            lcout => \generator_inst1.REGSTATZ0Z_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2249\,
            ce => \N__2195\,
            sr => \N__2145\
        );

    \generator_inst1.REGSTAT_34_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2366\,
            in2 => \_gnd_net_\,
            in3 => \N__1643\,
            lcout => \generator_inst1.REGSTATZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2249\,
            ce => \N__2195\,
            sr => \N__2145\
        );

    \generator_inst1.REGSTAT_37_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2369\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1655\,
            lcout => \generator_inst1.REGSTATZ0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2249\,
            ce => \N__2195\,
            sr => \N__2145\
        );

    \generator_inst1.REGSTAT_35_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2367\,
            in2 => \_gnd_net_\,
            in3 => \N__1667\,
            lcout => \generator_inst1.REGSTATZ0Z_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2249\,
            ce => \N__2195\,
            sr => \N__2145\
        );

    \generator_inst1.REGSTAT_36_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2368\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1661\,
            lcout => \generator_inst1.REGSTATZ0Z_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2249\,
            ce => \N__2195\,
            sr => \N__2145\
        );

    \generator_inst1.REGSTAT_39_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2371\,
            in2 => \_gnd_net_\,
            in3 => \N__1631\,
            lcout => \generator_inst1.REGSTATZ0Z_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2249\,
            ce => \N__2195\,
            sr => \N__2145\
        );

    \generator_inst1.REGSTAT_33_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2365\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1649\,
            lcout => \generator_inst1.REGSTATZ0Z_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2249\,
            ce => \N__2195\,
            sr => \N__2145\
        );

    \generator_inst1.REGSTAT_38_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2370\,
            in2 => \_gnd_net_\,
            in3 => \N__1637\,
            lcout => \generator_inst1.REGSTATZ0Z_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2249\,
            ce => \N__2195\,
            sr => \N__2145\
        );

    \generator_inst1.REGSTAT_41_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2323\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1826\,
            lcout => \generator_inst1.REGSTATZ0Z_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2248\,
            ce => \N__2194\,
            sr => \N__2143\
        );

    \generator_inst1.REGSTAT_40_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2322\,
            in2 => \_gnd_net_\,
            in3 => \N__1625\,
            lcout => \generator_inst1.REGSTATZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2248\,
            ce => \N__2194\,
            sr => \N__2143\
        );

    \generator_inst1.REGSTAT_44_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2326\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1808\,
            lcout => \generator_inst1.REGSTATZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2248\,
            ce => \N__2194\,
            sr => \N__2143\
        );

    \generator_inst1.REGSTAT_42_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2324\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1820\,
            lcout => \generator_inst1.REGSTATZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2248\,
            ce => \N__2194\,
            sr => \N__2143\
        );

    \generator_inst1.REGSTAT_43_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2325\,
            in2 => \_gnd_net_\,
            in3 => \N__1814\,
            lcout => \generator_inst1.REGSTATZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2248\,
            ce => \N__2194\,
            sr => \N__2143\
        );

    \generator_inst1.REGSTAT_45_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2327\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1802\,
            lcout => \generator_inst1.REGSTATZ0Z_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2248\,
            ce => \N__2194\,
            sr => \N__2143\
        );

    \SELDYN_ibuf_RNIKHL3_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1796\,
            lcout => \SELDYN_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RST_N_ibuf_RNIBJGC_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1706\,
            lcout => \RST_N_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.REGSTAT_80_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2607\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1880\,
            lcout => \generator_inst1.REGSTATZ0Z_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2261\,
            ce => \N__2206\,
            sr => \N__2156\
        );

    \generator_inst1.REGSTAT_82_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2609\,
            in2 => \_gnd_net_\,
            in3 => \N__1673\,
            lcout => \generator_inst1.REGSTATZ0Z_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2261\,
            ce => \N__2206\,
            sr => \N__2156\
        );

    \generator_inst1.REGSTAT_81_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2608\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1679\,
            lcout => \generator_inst1.REGSTATZ0Z_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2261\,
            ce => \N__2206\,
            sr => \N__2156\
        );

    \generator_inst1.REGSTAT_79_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2606\,
            in2 => \_gnd_net_\,
            in3 => \N__2018\,
            lcout => \generator_inst1.REGSTATZ0Z_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2261\,
            ce => \N__2206\,
            sr => \N__2156\
        );

    \generator_inst1.REGSTAT_83_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2610\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1874\,
            lcout => \generator_inst1.REGSTATZ0Z_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2261\,
            ce => \N__2206\,
            sr => \N__2156\
        );

    \generator_inst1.REGSTAT_2_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2586\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1904\,
            lcout => \generator_inst1.REGSTATZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2258\,
            ce => \N__2204\,
            sr => \N__2153\
        );

    \generator_inst1.REGSTAT_5_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2589\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1844\,
            lcout => \generator_inst1.REGSTATZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2258\,
            ce => \N__2204\,
            sr => \N__2153\
        );

    \generator_inst1.REGSTAT_3_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2587\,
            in2 => \_gnd_net_\,
            in3 => \N__1856\,
            lcout => \generator_inst1.REGSTATZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2258\,
            ce => \N__2204\,
            sr => \N__2153\
        );

    \generator_inst1.REGSTAT_4_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2588\,
            in2 => \_gnd_net_\,
            in3 => \N__1850\,
            lcout => \generator_inst1.REGSTATZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2258\,
            ce => \N__2204\,
            sr => \N__2153\
        );

    \generator_inst1.REGSTAT_25_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2578\,
            in2 => \_gnd_net_\,
            in3 => \N__1838\,
            lcout => \generator_inst1.REGSTATZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2255\,
            ce => \N__2201\,
            sr => \N__2150\
        );

    \generator_inst1.REGSTAT_24_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2577\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1832\,
            lcout => \generator_inst1.REGSTATZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2255\,
            ce => \N__2201\,
            sr => \N__2150\
        );

    \generator_inst1.REGSTAT_23_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2576\,
            in2 => \_gnd_net_\,
            in3 => \N__1928\,
            lcout => \generator_inst1.REGSTATZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2255\,
            ce => \N__2201\,
            sr => \N__2150\
        );

    \generator_inst1.REGSTAT_0_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2571\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \generator_inst1.REGSTATZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2255\,
            ce => \N__2201\,
            sr => \N__2150\
        );

    \generator_inst1.REGSTAT_20_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2573\,
            in2 => \_gnd_net_\,
            in3 => \N__1934\,
            lcout => \generator_inst1.REGSTATZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2255\,
            ce => \N__2201\,
            sr => \N__2150\
        );

    \generator_inst1.REGSTAT_22_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2575\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1916\,
            lcout => \generator_inst1.REGSTATZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2255\,
            ce => \N__2201\,
            sr => \N__2150\
        );

    \generator_inst1.REGSTAT_21_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2574\,
            in2 => \_gnd_net_\,
            in3 => \N__1922\,
            lcout => \generator_inst1.REGSTATZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2255\,
            ce => \N__2201\,
            sr => \N__2150\
        );

    \generator_inst1.REGSTAT_1_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2572\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1910\,
            lcout => \generator_inst1.REGSTATZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2255\,
            ce => \N__2201\,
            sr => \N__2150\
        );

    \generator_inst1.REGSTAT_30_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2569\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1886\,
            lcout => \generator_inst1.REGSTATZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2252\,
            ce => \N__2198\,
            sr => \N__2148\
        );

    \generator_inst1.REGSTAT_27_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2566\,
            in2 => \_gnd_net_\,
            in3 => \N__1988\,
            lcout => \generator_inst1.REGSTATZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2252\,
            ce => \N__2198\,
            sr => \N__2148\
        );

    \generator_inst1.REGSTAT_28_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2567\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1898\,
            lcout => \generator_inst1.REGSTATZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2252\,
            ce => \N__2198\,
            sr => \N__2148\
        );

    \generator_inst1.REGSTAT_29_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2568\,
            in2 => \_gnd_net_\,
            in3 => \N__1892\,
            lcout => \generator_inst1.REGSTATZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2252\,
            ce => \N__2198\,
            sr => \N__2148\
        );

    \generator_inst1.REGSTAT_26_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2565\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1994\,
            lcout => \generator_inst1.REGSTATZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2252\,
            ce => \N__2198\,
            sr => \N__2148\
        );

    \generator_inst1.REGSTAT_31_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2570\,
            in2 => \_gnd_net_\,
            in3 => \N__1982\,
            lcout => \generator_inst1.REGSTATZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2252\,
            ce => \N__2198\,
            sr => \N__2148\
        );

    \generator_inst1.REGSTAT_51_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2377\,
            in2 => \_gnd_net_\,
            in3 => \N__2036\,
            lcout => \generator_inst1.REGSTATZ0Z_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2250\,
            ce => \N__2196\,
            sr => \N__2144\
        );

    \generator_inst1.REGSTAT_47_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2373\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1952\,
            lcout => \generator_inst1.REGSTATZ0Z_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2250\,
            ce => \N__2196\,
            sr => \N__2144\
        );

    \generator_inst1.REGSTAT_53_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2379\,
            in2 => \_gnd_net_\,
            in3 => \N__1964\,
            lcout => \generator_inst1.REGSTATZ0Z_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2250\,
            ce => \N__2196\,
            sr => \N__2144\
        );

    \generator_inst1.REGSTAT_52_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2378\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1970\,
            lcout => \generator_inst1.REGSTATZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2250\,
            ce => \N__2196\,
            sr => \N__2144\
        );

    \generator_inst1.REGSTAT_46_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2372\,
            in2 => \_gnd_net_\,
            in3 => \N__1958\,
            lcout => \generator_inst1.REGSTATZ0Z_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2250\,
            ce => \N__2196\,
            sr => \N__2144\
        );

    \generator_inst1.REGSTAT_49_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2375\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1940\,
            lcout => \generator_inst1.REGSTATZ0Z_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2250\,
            ce => \N__2196\,
            sr => \N__2144\
        );

    \generator_inst1.REGSTAT_48_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2374\,
            in2 => \_gnd_net_\,
            in3 => \N__1946\,
            lcout => \generator_inst1.REGSTATZ0Z_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2250\,
            ce => \N__2196\,
            sr => \N__2144\
        );

    \generator_inst1.REGSTAT_50_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2376\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2042\,
            lcout => \generator_inst1.REGSTATZ0Z_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2250\,
            ce => \N__2196\,
            sr => \N__2144\
        );

    \generator_inst1.REGSTAT_76_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2599\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2012\,
            lcout => \generator_inst1.REGSTATZ0Z_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2262\,
            ce => \N__2207\,
            sr => \N__2157\
        );

    \generator_inst1.REGSTAT_77_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2600\,
            in2 => \_gnd_net_\,
            in3 => \N__2030\,
            lcout => \generator_inst1.REGSTATZ0Z_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2262\,
            ce => \N__2207\,
            sr => \N__2157\
        );

    \generator_inst1.REGSTAT_78_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2601\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2024\,
            lcout => \generator_inst1.REGSTATZ0Z_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2262\,
            ce => \N__2207\,
            sr => \N__2157\
        );

    \generator_inst1.REGSTAT_75_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2598\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2006\,
            lcout => \generator_inst1.REGSTATZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2262\,
            ce => \N__2207\,
            sr => \N__2157\
        );

    \generator_inst1.REGSTAT_74_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2597\,
            in2 => \_gnd_net_\,
            in3 => \N__2000\,
            lcout => \generator_inst1.REGSTATZ0Z_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2262\,
            ce => \N__2207\,
            sr => \N__2157\
        );

    \generator_inst1.REGSTAT_68_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2591\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2102\,
            lcout => \generator_inst1.REGSTATZ0Z_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2259\,
            ce => \N__2205\,
            sr => \N__2154\
        );

    \generator_inst1.REGSTAT_71_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2594\,
            in2 => \_gnd_net_\,
            in3 => \N__2096\,
            lcout => \generator_inst1.REGSTATZ0Z_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2259\,
            ce => \N__2205\,
            sr => \N__2154\
        );

    \generator_inst1.REGSTAT_73_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2596\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2072\,
            lcout => \generator_inst1.REGSTATZ0Z_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2259\,
            ce => \N__2205\,
            sr => \N__2154\
        );

    \generator_inst1.REGSTAT_67_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2590\,
            in2 => \_gnd_net_\,
            in3 => \N__2660\,
            lcout => \generator_inst1.REGSTATZ0Z_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2259\,
            ce => \N__2205\,
            sr => \N__2154\
        );

    \generator_inst1.REGSTAT_70_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2593\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2084\,
            lcout => \generator_inst1.REGSTATZ0Z_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2259\,
            ce => \N__2205\,
            sr => \N__2154\
        );

    \generator_inst1.REGSTAT_69_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2592\,
            in2 => \_gnd_net_\,
            in3 => \N__2090\,
            lcout => \generator_inst1.REGSTATZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2259\,
            ce => \N__2205\,
            sr => \N__2154\
        );

    \generator_inst1.REGSTAT_72_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2595\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2078\,
            lcout => \generator_inst1.REGSTATZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2259\,
            ce => \N__2205\,
            sr => \N__2154\
        );

    \generator_inst1.REGSTAT_64_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2583\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2066\,
            lcout => \generator_inst1.REGSTATZ0Z_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2256\,
            ce => \N__2202\,
            sr => \N__2151\
        );

    \generator_inst1.REGSTAT_60_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2579\,
            in2 => \_gnd_net_\,
            in3 => \N__2630\,
            lcout => \generator_inst1.REGSTATZ0Z_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2256\,
            ce => \N__2202\,
            sr => \N__2151\
        );

    \generator_inst1.REGSTAT_63_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2582\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2060\,
            lcout => \generator_inst1.REGSTATZ0Z_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2256\,
            ce => \N__2202\,
            sr => \N__2151\
        );

    \generator_inst1.REGSTAT_62_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2581\,
            in2 => \_gnd_net_\,
            in3 => \N__2048\,
            lcout => \generator_inst1.REGSTATZ0Z_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2256\,
            ce => \N__2202\,
            sr => \N__2151\
        );

    \generator_inst1.REGSTAT_61_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2580\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2054\,
            lcout => \generator_inst1.REGSTATZ0Z_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2256\,
            ce => \N__2202\,
            sr => \N__2151\
        );

    \generator_inst1.REGSTAT_66_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2585\,
            in2 => \_gnd_net_\,
            in3 => \N__2648\,
            lcout => \generator_inst1.REGSTATZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2256\,
            ce => \N__2202\,
            sr => \N__2151\
        );

    \generator_inst1.REGSTAT_65_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2584\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2654\,
            lcout => \generator_inst1.REGSTATZ0Z_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2256\,
            ce => \N__2202\,
            sr => \N__2151\
        );

    \generator_inst1.REGSTAT_57_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2383\,
            in2 => \_gnd_net_\,
            in3 => \N__2270\,
            lcout => \generator_inst1.REGSTATZ0Z_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2253\,
            ce => \N__2199\,
            sr => \N__2146\
        );

    \generator_inst1.REGSTAT_55_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2381\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2618\,
            lcout => \generator_inst1.REGSTATZ0Z_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2253\,
            ce => \N__2199\,
            sr => \N__2146\
        );

    \generator_inst1.REGSTAT_58_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2384\,
            in2 => \_gnd_net_\,
            in3 => \N__2642\,
            lcout => \generator_inst1.REGSTATZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2253\,
            ce => \N__2199\,
            sr => \N__2146\
        );

    \generator_inst1.REGSTAT_59_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2385\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2636\,
            lcout => \generator_inst1.REGSTATZ0Z_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2253\,
            ce => \N__2199\,
            sr => \N__2146\
        );

    \generator_inst1.REGSTAT_54_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2380\,
            in2 => \_gnd_net_\,
            in3 => \N__2624\,
            lcout => \generator_inst1.REGSTATZ0Z_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2253\,
            ce => \N__2199\,
            sr => \N__2146\
        );

    \generator_inst1.REGSTAT_56_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2382\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2276\,
            lcout => \generator_inst1.REGSTATZ0Z_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2253\,
            ce => \N__2199\,
            sr => \N__2146\
        );
end \INTERFACE\;
