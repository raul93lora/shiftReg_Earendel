// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 18 2025 09:13:17

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    generated_signal,
    RST_N,
    ENdin,
    CLK);

    output generated_signal;
    input RST_N;
    output ENdin;
    input CLK;

    wire N__1628;
    wire N__1627;
    wire N__1626;
    wire N__1617;
    wire N__1616;
    wire N__1615;
    wire N__1608;
    wire N__1607;
    wire N__1606;
    wire N__1599;
    wire N__1598;
    wire N__1597;
    wire N__1580;
    wire N__1579;
    wire N__1578;
    wire N__1575;
    wire N__1572;
    wire N__1569;
    wire N__1564;
    wire N__1561;
    wire N__1556;
    wire N__1553;
    wire N__1552;
    wire N__1551;
    wire N__1548;
    wire N__1545;
    wire N__1542;
    wire N__1535;
    wire N__1532;
    wire N__1531;
    wire N__1528;
    wire N__1525;
    wire N__1520;
    wire N__1517;
    wire N__1516;
    wire N__1515;
    wire N__1512;
    wire N__1507;
    wire N__1504;
    wire N__1499;
    wire N__1496;
    wire N__1495;
    wire N__1492;
    wire N__1489;
    wire N__1484;
    wire N__1481;
    wire N__1478;
    wire N__1477;
    wire N__1474;
    wire N__1471;
    wire N__1468;
    wire N__1463;
    wire N__1460;
    wire N__1459;
    wire N__1458;
    wire N__1457;
    wire N__1456;
    wire N__1455;
    wire N__1454;
    wire N__1453;
    wire N__1444;
    wire N__1435;
    wire N__1430;
    wire N__1427;
    wire N__1426;
    wire N__1423;
    wire N__1420;
    wire N__1415;
    wire N__1414;
    wire N__1413;
    wire N__1412;
    wire N__1411;
    wire N__1410;
    wire N__1409;
    wire N__1408;
    wire N__1407;
    wire N__1406;
    wire N__1405;
    wire N__1404;
    wire N__1379;
    wire N__1376;
    wire N__1373;
    wire N__1372;
    wire N__1371;
    wire N__1370;
    wire N__1369;
    wire N__1368;
    wire N__1367;
    wire N__1366;
    wire N__1365;
    wire N__1346;
    wire N__1343;
    wire N__1340;
    wire N__1339;
    wire N__1336;
    wire N__1333;
    wire N__1328;
    wire N__1325;
    wire N__1322;
    wire N__1319;
    wire N__1316;
    wire N__1315;
    wire N__1314;
    wire N__1313;
    wire N__1312;
    wire N__1311;
    wire N__1310;
    wire N__1309;
    wire N__1308;
    wire N__1307;
    wire N__1306;
    wire N__1305;
    wire N__1304;
    wire N__1303;
    wire N__1302;
    wire N__1299;
    wire N__1286;
    wire N__1269;
    wire N__1262;
    wire N__1261;
    wire N__1260;
    wire N__1259;
    wire N__1256;
    wire N__1253;
    wire N__1248;
    wire N__1241;
    wire N__1240;
    wire N__1235;
    wire N__1232;
    wire N__1229;
    wire N__1226;
    wire N__1225;
    wire N__1222;
    wire N__1219;
    wire N__1216;
    wire N__1211;
    wire N__1208;
    wire N__1205;
    wire N__1202;
    wire N__1199;
    wire N__1196;
    wire N__1193;
    wire N__1190;
    wire N__1187;
    wire N__1184;
    wire N__1181;
    wire N__1180;
    wire N__1179;
    wire N__1174;
    wire N__1171;
    wire N__1166;
    wire N__1163;
    wire N__1160;
    wire N__1157;
    wire N__1154;
    wire N__1151;
    wire N__1148;
    wire N__1145;
    wire N__1142;
    wire N__1139;
    wire N__1136;
    wire N__1133;
    wire N__1130;
    wire N__1127;
    wire N__1124;
    wire N__1121;
    wire N__1118;
    wire N__1115;
    wire N__1112;
    wire N__1109;
    wire N__1106;
    wire N__1103;
    wire N__1100;
    wire N__1097;
    wire N__1094;
    wire N__1091;
    wire N__1090;
    wire N__1087;
    wire N__1084;
    wire N__1079;
    wire N__1078;
    wire N__1077;
    wire N__1076;
    wire N__1073;
    wire N__1072;
    wire N__1071;
    wire N__1070;
    wire N__1061;
    wire N__1058;
    wire N__1053;
    wire N__1046;
    wire N__1045;
    wire N__1044;
    wire N__1043;
    wire N__1040;
    wire N__1035;
    wire N__1032;
    wire N__1025;
    wire N__1022;
    wire N__1019;
    wire N__1016;
    wire N__1013;
    wire N__1010;
    wire N__1007;
    wire N__1004;
    wire N__1001;
    wire N__998;
    wire N__995;
    wire N__994;
    wire N__993;
    wire N__990;
    wire N__989;
    wire N__988;
    wire N__985;
    wire N__984;
    wire N__981;
    wire N__974;
    wire N__969;
    wire N__962;
    wire N__959;
    wire N__956;
    wire N__955;
    wire N__952;
    wire N__951;
    wire N__950;
    wire N__949;
    wire N__948;
    wire N__947;
    wire N__946;
    wire N__945;
    wire N__942;
    wire N__939;
    wire N__936;
    wire N__929;
    wire N__922;
    wire N__911;
    wire N__908;
    wire N__905;
    wire N__902;
    wire N__899;
    wire N__896;
    wire N__893;
    wire N__892;
    wire N__889;
    wire N__886;
    wire N__881;
    wire N__878;
    wire N__877;
    wire N__876;
    wire N__875;
    wire N__874;
    wire N__869;
    wire N__862;
    wire N__857;
    wire N__856;
    wire N__855;
    wire N__854;
    wire N__851;
    wire N__848;
    wire N__843;
    wire N__840;
    wire N__833;
    wire N__832;
    wire N__829;
    wire N__828;
    wire N__821;
    wire N__818;
    wire N__815;
    wire N__812;
    wire N__809;
    wire N__808;
    wire N__807;
    wire N__804;
    wire N__799;
    wire N__796;
    wire N__793;
    wire N__788;
    wire N__785;
    wire N__782;
    wire N__779;
    wire N__776;
    wire N__773;
    wire N__770;
    wire N__769;
    wire N__768;
    wire N__767;
    wire N__766;
    wire N__755;
    wire N__752;
    wire N__751;
    wire N__750;
    wire N__749;
    wire N__746;
    wire N__739;
    wire N__734;
    wire N__731;
    wire N__730;
    wire N__729;
    wire N__728;
    wire N__725;
    wire N__722;
    wire N__719;
    wire N__718;
    wire N__715;
    wire N__706;
    wire VCCG0;
    wire GNDG0;
    wire RST_N_c_i;
    wire \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_ ;
    wire \fsm_shiftRegs_inst1.counterZ0Z_0 ;
    wire \fsm_shiftRegs_inst1.counterZ0Z_1 ;
    wire \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3_cascade_ ;
    wire \fsm_shiftRegs_inst1.counterZ0Z_3 ;
    wire \fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_ ;
    wire \fsm_shiftRegs_inst1.N_123_1 ;
    wire \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_ ;
    wire \fsm_shiftRegs_inst1.counterDYNZ0Z_1 ;
    wire \fsm_shiftRegs_inst1.counterDYNZ0Z_2 ;
    wire \fsm_shiftRegs_inst1.counterDYNZ0Z_3 ;
    wire RST_N_c;
    wire \fsm_shiftRegs_inst1.current_stateZ0Z_1 ;
    wire \fsm_shiftRegs_inst1.counterZ0Z_2 ;
    wire \fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2 ;
    wire ENdin_c;
    wire \fsm_shiftRegs_inst1.counterDYNZ0Z_0 ;
    wire \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3 ;
    wire \fsm_shiftRegs_inst1.current_stateZ0Z_2 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_10 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_13 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_14 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_15 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_11 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_12 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_8 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_9 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_6 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_7 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_2 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_3 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_4 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_5 ;
    wire \fsm_shiftRegs_inst1.un1_current_state4_0 ;
    wire \fsm_shiftRegs_inst1.current_stateZ0Z_3 ;
    wire \fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_ ;
    wire \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_ ;
    wire \fsm_shiftRegs_inst1.current_stateZ0Z_0 ;
    wire \fsm_shiftRegs_inst1.current_stateZ0Z_4 ;
    wire \fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0 ;
    wire SELSTAT;
    wire signal_out_fsm;
    wire SELDYN;
    wire generated_signal_c;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_0 ;
    wire bfn_16_16_0_;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_1 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_0 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_2 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_1 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_3 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_2 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_4 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_3 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_5 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_4 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_6 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_5 ;
    wire \fsm_shiftRegs_inst1.current_state_i_4 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_6 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_7 ;
    wire _gnd_net_;
    wire CLK_c_g;
    wire RST_N_c_i_g;

    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__1626),
            .GLOBALBUFFEROUTPUT(CLK_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__1628),
            .DIN(N__1627),
            .DOUT(N__1626),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__1628),
            .PADOUT(N__1627),
            .PADIN(N__1626),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RST_N_ibuf_iopad (
            .OE(N__1617),
            .DIN(N__1616),
            .DOUT(N__1615),
            .PACKAGEPIN(RST_N));
    defparam RST_N_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RST_N_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RST_N_ibuf_preio (
            .PADOEN(N__1617),
            .PADOUT(N__1616),
            .PADIN(N__1615),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RST_N_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD generated_signal_obuf_iopad (
            .OE(N__1608),
            .DIN(N__1607),
            .DOUT(N__1606),
            .PACKAGEPIN(generated_signal));
    defparam generated_signal_obuf_preio.NEG_TRIGGER=1'b0;
    defparam generated_signal_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO generated_signal_obuf_preio (
            .PADOEN(N__1608),
            .PADOUT(N__1607),
            .PADIN(N__1606),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1205),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ENdin_obuf_iopad (
            .OE(N__1599),
            .DIN(N__1598),
            .DOUT(N__1597),
            .PACKAGEPIN(ENdin));
    defparam ENdin_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ENdin_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ENdin_obuf_preio (
            .PADOEN(N__1599),
            .PADOUT(N__1598),
            .PADIN(N__1597),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1016),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__354 (
            .O(N__1580),
            .I(N__1575));
    CascadeMux I__353 (
            .O(N__1579),
            .I(N__1572));
    CascadeMux I__352 (
            .O(N__1578),
            .I(N__1569));
    InMux I__351 (
            .O(N__1575),
            .I(N__1564));
    InMux I__350 (
            .O(N__1572),
            .I(N__1564));
    InMux I__349 (
            .O(N__1569),
            .I(N__1561));
    LocalMux I__348 (
            .O(N__1564),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_1 ));
    LocalMux I__347 (
            .O(N__1561),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_1 ));
    InMux I__346 (
            .O(N__1556),
            .I(\fsm_shiftRegs_inst1.counter2_cry_0 ));
    InMux I__345 (
            .O(N__1553),
            .I(N__1548));
    InMux I__344 (
            .O(N__1552),
            .I(N__1545));
    InMux I__343 (
            .O(N__1551),
            .I(N__1542));
    LocalMux I__342 (
            .O(N__1548),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_2 ));
    LocalMux I__341 (
            .O(N__1545),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_2 ));
    LocalMux I__340 (
            .O(N__1542),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_2 ));
    InMux I__339 (
            .O(N__1535),
            .I(\fsm_shiftRegs_inst1.counter2_cry_1 ));
    InMux I__338 (
            .O(N__1532),
            .I(N__1528));
    InMux I__337 (
            .O(N__1531),
            .I(N__1525));
    LocalMux I__336 (
            .O(N__1528),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_3 ));
    LocalMux I__335 (
            .O(N__1525),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_3 ));
    InMux I__334 (
            .O(N__1520),
            .I(\fsm_shiftRegs_inst1.counter2_cry_2 ));
    CascadeMux I__333 (
            .O(N__1517),
            .I(N__1512));
    InMux I__332 (
            .O(N__1516),
            .I(N__1507));
    InMux I__331 (
            .O(N__1515),
            .I(N__1507));
    InMux I__330 (
            .O(N__1512),
            .I(N__1504));
    LocalMux I__329 (
            .O(N__1507),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_4 ));
    LocalMux I__328 (
            .O(N__1504),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_4 ));
    InMux I__327 (
            .O(N__1499),
            .I(\fsm_shiftRegs_inst1.counter2_cry_3 ));
    InMux I__326 (
            .O(N__1496),
            .I(N__1492));
    InMux I__325 (
            .O(N__1495),
            .I(N__1489));
    LocalMux I__324 (
            .O(N__1492),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_5 ));
    LocalMux I__323 (
            .O(N__1489),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_5 ));
    InMux I__322 (
            .O(N__1484),
            .I(\fsm_shiftRegs_inst1.counter2_cry_4 ));
    CascadeMux I__321 (
            .O(N__1481),
            .I(N__1478));
    InMux I__320 (
            .O(N__1478),
            .I(N__1474));
    InMux I__319 (
            .O(N__1477),
            .I(N__1471));
    LocalMux I__318 (
            .O(N__1474),
            .I(N__1468));
    LocalMux I__317 (
            .O(N__1471),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_6 ));
    Odrv4 I__316 (
            .O(N__1468),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_6 ));
    InMux I__315 (
            .O(N__1463),
            .I(\fsm_shiftRegs_inst1.counter2_cry_5 ));
    InMux I__314 (
            .O(N__1460),
            .I(N__1444));
    InMux I__313 (
            .O(N__1459),
            .I(N__1444));
    InMux I__312 (
            .O(N__1458),
            .I(N__1444));
    InMux I__311 (
            .O(N__1457),
            .I(N__1444));
    InMux I__310 (
            .O(N__1456),
            .I(N__1435));
    InMux I__309 (
            .O(N__1455),
            .I(N__1435));
    InMux I__308 (
            .O(N__1454),
            .I(N__1435));
    InMux I__307 (
            .O(N__1453),
            .I(N__1435));
    LocalMux I__306 (
            .O(N__1444),
            .I(\fsm_shiftRegs_inst1.current_state_i_4 ));
    LocalMux I__305 (
            .O(N__1435),
            .I(\fsm_shiftRegs_inst1.current_state_i_4 ));
    InMux I__304 (
            .O(N__1430),
            .I(\fsm_shiftRegs_inst1.counter2_cry_6 ));
    InMux I__303 (
            .O(N__1427),
            .I(N__1423));
    InMux I__302 (
            .O(N__1426),
            .I(N__1420));
    LocalMux I__301 (
            .O(N__1423),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_7 ));
    LocalMux I__300 (
            .O(N__1420),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_7 ));
    ClkMux I__299 (
            .O(N__1415),
            .I(N__1379));
    ClkMux I__298 (
            .O(N__1414),
            .I(N__1379));
    ClkMux I__297 (
            .O(N__1413),
            .I(N__1379));
    ClkMux I__296 (
            .O(N__1412),
            .I(N__1379));
    ClkMux I__295 (
            .O(N__1411),
            .I(N__1379));
    ClkMux I__294 (
            .O(N__1410),
            .I(N__1379));
    ClkMux I__293 (
            .O(N__1409),
            .I(N__1379));
    ClkMux I__292 (
            .O(N__1408),
            .I(N__1379));
    ClkMux I__291 (
            .O(N__1407),
            .I(N__1379));
    ClkMux I__290 (
            .O(N__1406),
            .I(N__1379));
    ClkMux I__289 (
            .O(N__1405),
            .I(N__1379));
    ClkMux I__288 (
            .O(N__1404),
            .I(N__1379));
    GlobalMux I__287 (
            .O(N__1379),
            .I(N__1376));
    gio2CtrlBuf I__286 (
            .O(N__1376),
            .I(CLK_c_g));
    SRMux I__285 (
            .O(N__1373),
            .I(N__1346));
    SRMux I__284 (
            .O(N__1372),
            .I(N__1346));
    SRMux I__283 (
            .O(N__1371),
            .I(N__1346));
    SRMux I__282 (
            .O(N__1370),
            .I(N__1346));
    SRMux I__281 (
            .O(N__1369),
            .I(N__1346));
    SRMux I__280 (
            .O(N__1368),
            .I(N__1346));
    SRMux I__279 (
            .O(N__1367),
            .I(N__1346));
    SRMux I__278 (
            .O(N__1366),
            .I(N__1346));
    SRMux I__277 (
            .O(N__1365),
            .I(N__1346));
    GlobalMux I__276 (
            .O(N__1346),
            .I(N__1343));
    gio2CtrlBuf I__275 (
            .O(N__1343),
            .I(RST_N_c_i_g));
    InMux I__274 (
            .O(N__1340),
            .I(N__1336));
    InMux I__273 (
            .O(N__1339),
            .I(N__1333));
    LocalMux I__272 (
            .O(N__1336),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_3 ));
    LocalMux I__271 (
            .O(N__1333),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_3 ));
    CascadeMux I__270 (
            .O(N__1328),
            .I(\fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_ ));
    CascadeMux I__269 (
            .O(N__1325),
            .I(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_ ));
    CascadeMux I__268 (
            .O(N__1322),
            .I(N__1319));
    InMux I__267 (
            .O(N__1319),
            .I(N__1316));
    LocalMux I__266 (
            .O(N__1316),
            .I(N__1299));
    InMux I__265 (
            .O(N__1315),
            .I(N__1286));
    InMux I__264 (
            .O(N__1314),
            .I(N__1286));
    InMux I__263 (
            .O(N__1313),
            .I(N__1286));
    InMux I__262 (
            .O(N__1312),
            .I(N__1286));
    InMux I__261 (
            .O(N__1311),
            .I(N__1286));
    InMux I__260 (
            .O(N__1310),
            .I(N__1286));
    InMux I__259 (
            .O(N__1309),
            .I(N__1269));
    InMux I__258 (
            .O(N__1308),
            .I(N__1269));
    InMux I__257 (
            .O(N__1307),
            .I(N__1269));
    InMux I__256 (
            .O(N__1306),
            .I(N__1269));
    InMux I__255 (
            .O(N__1305),
            .I(N__1269));
    InMux I__254 (
            .O(N__1304),
            .I(N__1269));
    InMux I__253 (
            .O(N__1303),
            .I(N__1269));
    InMux I__252 (
            .O(N__1302),
            .I(N__1269));
    Odrv12 I__251 (
            .O(N__1299),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_0 ));
    LocalMux I__250 (
            .O(N__1286),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_0 ));
    LocalMux I__249 (
            .O(N__1269),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_0 ));
    InMux I__248 (
            .O(N__1262),
            .I(N__1256));
    InMux I__247 (
            .O(N__1261),
            .I(N__1253));
    InMux I__246 (
            .O(N__1260),
            .I(N__1248));
    InMux I__245 (
            .O(N__1259),
            .I(N__1248));
    LocalMux I__244 (
            .O(N__1256),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_4 ));
    LocalMux I__243 (
            .O(N__1253),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_4 ));
    LocalMux I__242 (
            .O(N__1248),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_4 ));
    InMux I__241 (
            .O(N__1241),
            .I(N__1235));
    InMux I__240 (
            .O(N__1240),
            .I(N__1235));
    LocalMux I__239 (
            .O(N__1235),
            .I(\fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0 ));
    InMux I__238 (
            .O(N__1232),
            .I(N__1229));
    LocalMux I__237 (
            .O(N__1229),
            .I(SELSTAT));
    InMux I__236 (
            .O(N__1226),
            .I(N__1222));
    InMux I__235 (
            .O(N__1225),
            .I(N__1219));
    LocalMux I__234 (
            .O(N__1222),
            .I(N__1216));
    LocalMux I__233 (
            .O(N__1219),
            .I(signal_out_fsm));
    Odrv12 I__232 (
            .O(N__1216),
            .I(signal_out_fsm));
    InMux I__231 (
            .O(N__1211),
            .I(N__1208));
    LocalMux I__230 (
            .O(N__1208),
            .I(SELDYN));
    IoInMux I__229 (
            .O(N__1205),
            .I(N__1202));
    LocalMux I__228 (
            .O(N__1202),
            .I(N__1199));
    IoSpan4Mux I__227 (
            .O(N__1199),
            .I(N__1196));
    IoSpan4Mux I__226 (
            .O(N__1196),
            .I(N__1193));
    Sp12to4 I__225 (
            .O(N__1193),
            .I(N__1190));
    Span12Mux_s7_h I__224 (
            .O(N__1190),
            .I(N__1187));
    Span12Mux_v I__223 (
            .O(N__1187),
            .I(N__1184));
    Odrv12 I__222 (
            .O(N__1184),
            .I(generated_signal_c));
    InMux I__221 (
            .O(N__1181),
            .I(N__1174));
    InMux I__220 (
            .O(N__1180),
            .I(N__1174));
    InMux I__219 (
            .O(N__1179),
            .I(N__1171));
    LocalMux I__218 (
            .O(N__1174),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_0 ));
    LocalMux I__217 (
            .O(N__1171),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_0 ));
    InMux I__216 (
            .O(N__1166),
            .I(bfn_16_16_0_));
    InMux I__215 (
            .O(N__1163),
            .I(N__1160));
    LocalMux I__214 (
            .O(N__1160),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_14 ));
    InMux I__213 (
            .O(N__1157),
            .I(N__1154));
    LocalMux I__212 (
            .O(N__1154),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_15 ));
    InMux I__211 (
            .O(N__1151),
            .I(N__1148));
    LocalMux I__210 (
            .O(N__1148),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_11 ));
    InMux I__209 (
            .O(N__1145),
            .I(N__1142));
    LocalMux I__208 (
            .O(N__1142),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_12 ));
    InMux I__207 (
            .O(N__1139),
            .I(N__1136));
    LocalMux I__206 (
            .O(N__1136),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_8 ));
    InMux I__205 (
            .O(N__1133),
            .I(N__1130));
    LocalMux I__204 (
            .O(N__1130),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_9 ));
    InMux I__203 (
            .O(N__1127),
            .I(N__1124));
    LocalMux I__202 (
            .O(N__1124),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_6 ));
    InMux I__201 (
            .O(N__1121),
            .I(N__1118));
    LocalMux I__200 (
            .O(N__1118),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_7 ));
    InMux I__199 (
            .O(N__1115),
            .I(N__1112));
    LocalMux I__198 (
            .O(N__1112),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_2 ));
    InMux I__197 (
            .O(N__1109),
            .I(N__1106));
    LocalMux I__196 (
            .O(N__1106),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_3 ));
    InMux I__195 (
            .O(N__1103),
            .I(N__1100));
    LocalMux I__194 (
            .O(N__1100),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_4 ));
    InMux I__193 (
            .O(N__1097),
            .I(N__1094));
    LocalMux I__192 (
            .O(N__1094),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_5 ));
    CEMux I__191 (
            .O(N__1091),
            .I(N__1087));
    CEMux I__190 (
            .O(N__1090),
            .I(N__1084));
    LocalMux I__189 (
            .O(N__1087),
            .I(\fsm_shiftRegs_inst1.un1_current_state4_0 ));
    LocalMux I__188 (
            .O(N__1084),
            .I(\fsm_shiftRegs_inst1.un1_current_state4_0 ));
    CascadeMux I__187 (
            .O(N__1079),
            .I(N__1073));
    InMux I__186 (
            .O(N__1078),
            .I(N__1061));
    InMux I__185 (
            .O(N__1077),
            .I(N__1061));
    InMux I__184 (
            .O(N__1076),
            .I(N__1061));
    InMux I__183 (
            .O(N__1073),
            .I(N__1061));
    InMux I__182 (
            .O(N__1072),
            .I(N__1058));
    InMux I__181 (
            .O(N__1071),
            .I(N__1053));
    InMux I__180 (
            .O(N__1070),
            .I(N__1053));
    LocalMux I__179 (
            .O(N__1061),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_1 ));
    LocalMux I__178 (
            .O(N__1058),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_1 ));
    LocalMux I__177 (
            .O(N__1053),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_1 ));
    InMux I__176 (
            .O(N__1046),
            .I(N__1040));
    InMux I__175 (
            .O(N__1045),
            .I(N__1035));
    InMux I__174 (
            .O(N__1044),
            .I(N__1035));
    InMux I__173 (
            .O(N__1043),
            .I(N__1032));
    LocalMux I__172 (
            .O(N__1040),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_2 ));
    LocalMux I__171 (
            .O(N__1035),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_2 ));
    LocalMux I__170 (
            .O(N__1032),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_2 ));
    InMux I__169 (
            .O(N__1025),
            .I(N__1022));
    LocalMux I__168 (
            .O(N__1022),
            .I(N__1019));
    Odrv4 I__167 (
            .O(N__1019),
            .I(\fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2 ));
    IoInMux I__166 (
            .O(N__1016),
            .I(N__1013));
    LocalMux I__165 (
            .O(N__1013),
            .I(N__1010));
    IoSpan4Mux I__164 (
            .O(N__1010),
            .I(N__1007));
    Span4Mux_s3_h I__163 (
            .O(N__1007),
            .I(N__1004));
    Sp12to4 I__162 (
            .O(N__1004),
            .I(N__1001));
    Span12Mux_h I__161 (
            .O(N__1001),
            .I(N__998));
    Odrv12 I__160 (
            .O(N__998),
            .I(ENdin_c));
    CascadeMux I__159 (
            .O(N__995),
            .I(N__990));
    CascadeMux I__158 (
            .O(N__994),
            .I(N__985));
    InMux I__157 (
            .O(N__993),
            .I(N__981));
    InMux I__156 (
            .O(N__990),
            .I(N__974));
    InMux I__155 (
            .O(N__989),
            .I(N__974));
    InMux I__154 (
            .O(N__988),
            .I(N__974));
    InMux I__153 (
            .O(N__985),
            .I(N__969));
    InMux I__152 (
            .O(N__984),
            .I(N__969));
    LocalMux I__151 (
            .O(N__981),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_0 ));
    LocalMux I__150 (
            .O(N__974),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_0 ));
    LocalMux I__149 (
            .O(N__969),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_0 ));
    InMux I__148 (
            .O(N__962),
            .I(N__959));
    LocalMux I__147 (
            .O(N__959),
            .I(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3 ));
    CascadeMux I__146 (
            .O(N__956),
            .I(N__952));
    InMux I__145 (
            .O(N__955),
            .I(N__942));
    InMux I__144 (
            .O(N__952),
            .I(N__939));
    InMux I__143 (
            .O(N__951),
            .I(N__936));
    InMux I__142 (
            .O(N__950),
            .I(N__929));
    InMux I__141 (
            .O(N__949),
            .I(N__929));
    InMux I__140 (
            .O(N__948),
            .I(N__929));
    InMux I__139 (
            .O(N__947),
            .I(N__922));
    InMux I__138 (
            .O(N__946),
            .I(N__922));
    InMux I__137 (
            .O(N__945),
            .I(N__922));
    LocalMux I__136 (
            .O(N__942),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ));
    LocalMux I__135 (
            .O(N__939),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ));
    LocalMux I__134 (
            .O(N__936),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ));
    LocalMux I__133 (
            .O(N__929),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ));
    LocalMux I__132 (
            .O(N__922),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ));
    InMux I__131 (
            .O(N__911),
            .I(N__908));
    LocalMux I__130 (
            .O(N__908),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_10 ));
    InMux I__129 (
            .O(N__905),
            .I(N__902));
    LocalMux I__128 (
            .O(N__902),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_13 ));
    CascadeMux I__127 (
            .O(N__899),
            .I(\fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_ ));
    InMux I__126 (
            .O(N__896),
            .I(N__893));
    LocalMux I__125 (
            .O(N__893),
            .I(N__889));
    InMux I__124 (
            .O(N__892),
            .I(N__886));
    Odrv4 I__123 (
            .O(N__889),
            .I(\fsm_shiftRegs_inst1.N_123_1 ));
    LocalMux I__122 (
            .O(N__886),
            .I(\fsm_shiftRegs_inst1.N_123_1 ));
    CascadeMux I__121 (
            .O(N__881),
            .I(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_ ));
    InMux I__120 (
            .O(N__878),
            .I(N__869));
    InMux I__119 (
            .O(N__877),
            .I(N__869));
    InMux I__118 (
            .O(N__876),
            .I(N__862));
    InMux I__117 (
            .O(N__875),
            .I(N__862));
    InMux I__116 (
            .O(N__874),
            .I(N__862));
    LocalMux I__115 (
            .O(N__869),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_1 ));
    LocalMux I__114 (
            .O(N__862),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_1 ));
    CascadeMux I__113 (
            .O(N__857),
            .I(N__851));
    InMux I__112 (
            .O(N__856),
            .I(N__848));
    InMux I__111 (
            .O(N__855),
            .I(N__843));
    InMux I__110 (
            .O(N__854),
            .I(N__843));
    InMux I__109 (
            .O(N__851),
            .I(N__840));
    LocalMux I__108 (
            .O(N__848),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_2 ));
    LocalMux I__107 (
            .O(N__843),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_2 ));
    LocalMux I__106 (
            .O(N__840),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_2 ));
    CascadeMux I__105 (
            .O(N__833),
            .I(N__829));
    InMux I__104 (
            .O(N__832),
            .I(N__821));
    InMux I__103 (
            .O(N__829),
            .I(N__821));
    InMux I__102 (
            .O(N__828),
            .I(N__821));
    LocalMux I__101 (
            .O(N__821),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_3 ));
    InMux I__100 (
            .O(N__818),
            .I(N__815));
    LocalMux I__99 (
            .O(N__815),
            .I(N__812));
    Span4Mux_v I__98 (
            .O(N__812),
            .I(N__809));
    Span4Mux_v I__97 (
            .O(N__809),
            .I(N__804));
    InMux I__96 (
            .O(N__808),
            .I(N__799));
    InMux I__95 (
            .O(N__807),
            .I(N__799));
    Sp12to4 I__94 (
            .O(N__804),
            .I(N__796));
    LocalMux I__93 (
            .O(N__799),
            .I(N__793));
    Span12Mux_h I__92 (
            .O(N__796),
            .I(N__788));
    Span12Mux_v I__91 (
            .O(N__793),
            .I(N__788));
    Span12Mux_h I__90 (
            .O(N__788),
            .I(N__785));
    Odrv12 I__89 (
            .O(N__785),
            .I(RST_N_c));
    IoInMux I__88 (
            .O(N__782),
            .I(N__779));
    LocalMux I__87 (
            .O(N__779),
            .I(N__776));
    Odrv12 I__86 (
            .O(N__776),
            .I(RST_N_c_i));
    CascadeMux I__85 (
            .O(N__773),
            .I(\fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_ ));
    InMux I__84 (
            .O(N__770),
            .I(N__755));
    InMux I__83 (
            .O(N__769),
            .I(N__755));
    InMux I__82 (
            .O(N__768),
            .I(N__755));
    InMux I__81 (
            .O(N__767),
            .I(N__755));
    InMux I__80 (
            .O(N__766),
            .I(N__755));
    LocalMux I__79 (
            .O(N__755),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_0 ));
    InMux I__78 (
            .O(N__752),
            .I(N__746));
    InMux I__77 (
            .O(N__751),
            .I(N__739));
    InMux I__76 (
            .O(N__750),
            .I(N__739));
    InMux I__75 (
            .O(N__749),
            .I(N__739));
    LocalMux I__74 (
            .O(N__746),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_1 ));
    LocalMux I__73 (
            .O(N__739),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_1 ));
    CascadeMux I__72 (
            .O(N__734),
            .I(\fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3_cascade_ ));
    CascadeMux I__71 (
            .O(N__731),
            .I(N__725));
    CascadeMux I__70 (
            .O(N__730),
            .I(N__722));
    CascadeMux I__69 (
            .O(N__729),
            .I(N__719));
    InMux I__68 (
            .O(N__728),
            .I(N__715));
    InMux I__67 (
            .O(N__725),
            .I(N__706));
    InMux I__66 (
            .O(N__722),
            .I(N__706));
    InMux I__65 (
            .O(N__719),
            .I(N__706));
    InMux I__64 (
            .O(N__718),
            .I(N__706));
    LocalMux I__63 (
            .O(N__715),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_3 ));
    LocalMux I__62 (
            .O(N__706),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_3 ));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_16_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB RST_N_ibuf_RNIBJGC_0 (
            .USERSIGNALTOGLOBALBUFFER(N__782),
            .GLOBALBUFFEROUTPUT(RST_N_c_i_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam RST_N_ibuf_RNIBJGC_LC_4_16_1.C_ON=1'b0;
    defparam RST_N_ibuf_RNIBJGC_LC_4_16_1.SEQ_MODE=4'b0000;
    defparam RST_N_ibuf_RNIBJGC_LC_4_16_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 RST_N_ibuf_RNIBJGC_LC_4_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__818),
            .lcout(RST_N_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_2_LC_13_14_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_2_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_2_LC_13_14_0 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \fsm_shiftRegs_inst1.counter_RNO_0_2_LC_13_14_0  (
            .in0(N__767),
            .in1(N__750),
            .in2(N__729),
            .in3(N__1044),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counter_2_LC_13_14_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_2_LC_13_14_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter_2_LC_13_14_1 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \fsm_shiftRegs_inst1.counter_2_LC_13_14_1  (
            .in0(N__1076),
            .in1(_gnd_net_),
            .in2(N__773),
            .in3(_gnd_net_),
            .lcout(\fsm_shiftRegs_inst1.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1405),
            .ce(),
            .sr(N__1366));
    defparam \fsm_shiftRegs_inst1.counter_0_LC_13_14_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_0_LC_13_14_2 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter_0_LC_13_14_2 .LUT_INIT=16'b1010010100000000;
    LogicCell40 \fsm_shiftRegs_inst1.counter_0_LC_13_14_2  (
            .in0(N__769),
            .in1(_gnd_net_),
            .in2(N__731),
            .in3(N__1078),
            .lcout(\fsm_shiftRegs_inst1.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1405),
            .ce(),
            .sr(N__1366));
    defparam \fsm_shiftRegs_inst1.counter_RNIC589_1_LC_13_14_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_RNIC589_1_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.counter_RNIC589_1_LC_13_14_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \fsm_shiftRegs_inst1.counter_RNIC589_1_LC_13_14_3  (
            .in0(N__749),
            .in1(N__766),
            .in2(_gnd_net_),
            .in3(N__718),
            .lcout(\fsm_shiftRegs_inst1.N_123_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counter_1_LC_13_14_5 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_1_LC_13_14_5 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter_1_LC_13_14_5 .LUT_INIT=16'b1001000011000000;
    LogicCell40 \fsm_shiftRegs_inst1.counter_1_LC_13_14_5  (
            .in0(N__728),
            .in1(N__752),
            .in2(N__1079),
            .in3(N__770),
            .lcout(\fsm_shiftRegs_inst1.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1405),
            .ce(),
            .sr(N__1366));
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_3_LC_13_14_6 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_3_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_3_LC_13_14_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \fsm_shiftRegs_inst1.counter_RNO_0_3_LC_13_14_6  (
            .in0(N__768),
            .in1(N__751),
            .in2(N__730),
            .in3(N__1045),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counter_3_LC_13_14_7 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_3_LC_13_14_7 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter_3_LC_13_14_7 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \fsm_shiftRegs_inst1.counter_3_LC_13_14_7  (
            .in0(N__1077),
            .in1(_gnd_net_),
            .in2(N__734),
            .in3(_gnd_net_),
            .lcout(\fsm_shiftRegs_inst1.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1405),
            .ce(),
            .sr(N__1366));
    defparam \fsm_shiftRegs_inst1.current_state_1_LC_13_15_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_1_LC_13_15_3 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.current_state_1_LC_13_15_3 .LUT_INIT=16'b1111100011111010;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_1_LC_13_15_3  (
            .in0(N__1072),
            .in1(N__1046),
            .in2(N__1322),
            .in3(N__892),
            .lcout(\fsm_shiftRegs_inst1.current_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1404),
            .ce(),
            .sr(N__1365));
    defparam \fsm_shiftRegs_inst1.counterDYN_1_LC_14_13_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counterDYN_1_LC_14_13_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counterDYN_1_LC_14_13_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \fsm_shiftRegs_inst1.counterDYN_1_LC_14_13_1  (
            .in0(N__948),
            .in1(N__989),
            .in2(_gnd_net_),
            .in3(N__878),
            .lcout(\fsm_shiftRegs_inst1.counterDYNZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1411),
            .ce(),
            .sr(N__1369));
    defparam \fsm_shiftRegs_inst1.counterDYN_2_LC_14_13_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counterDYN_2_LC_14_13_2 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counterDYN_2_LC_14_13_2 .LUT_INIT=16'b0100110010000000;
    LogicCell40 \fsm_shiftRegs_inst1.counterDYN_2_LC_14_13_2  (
            .in0(N__877),
            .in1(N__950),
            .in2(N__995),
            .in3(N__856),
            .lcout(\fsm_shiftRegs_inst1.counterDYNZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1411),
            .ce(),
            .sr(N__1369));
    defparam \fsm_shiftRegs_inst1.counterDYN_0_LC_14_13_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counterDYN_0_LC_14_13_3 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counterDYN_0_LC_14_13_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \fsm_shiftRegs_inst1.counterDYN_0_LC_14_13_3  (
            .in0(N__949),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__988),
            .lcout(\fsm_shiftRegs_inst1.counterDYNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1411),
            .ce(),
            .sr(N__1369));
    defparam \fsm_shiftRegs_inst1.counterDYN_RNO_0_3_LC_14_14_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counterDYN_RNO_0_3_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.counterDYN_RNO_0_3_LC_14_14_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \fsm_shiftRegs_inst1.counterDYN_RNO_0_3_LC_14_14_0  (
            .in0(N__854),
            .in1(N__875),
            .in2(N__833),
            .in3(N__984),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counterDYN_3_LC_14_14_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counterDYN_3_LC_14_14_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counterDYN_3_LC_14_14_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fsm_shiftRegs_inst1.counterDYN_3_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__899),
            .in3(N__947),
            .lcout(\fsm_shiftRegs_inst1.counterDYNZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1408),
            .ce(),
            .sr(N__1368));
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_2_LC_14_14_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_2_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_2_LC_14_14_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNO_0_2_LC_14_14_3  (
            .in0(N__876),
            .in1(N__855),
            .in2(N__994),
            .in3(N__832),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_2_LC_14_14_4 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_2_LC_14_14_4 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.current_state_2_LC_14_14_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_2_LC_14_14_4  (
            .in0(N__946),
            .in1(N__896),
            .in2(N__881),
            .in3(N__1025),
            .lcout(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1408),
            .ce(),
            .sr(N__1368));
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_3_LC_14_14_5 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_3_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_3_LC_14_14_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNO_0_3_LC_14_14_5  (
            .in0(N__874),
            .in1(N__945),
            .in2(N__857),
            .in3(N__828),
            .lcout(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.signal_out_LC_14_15_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.signal_out_LC_14_15_0 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.signal_out_LC_14_15_0 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \fsm_shiftRegs_inst1.signal_out_LC_14_15_0  (
            .in0(N__1225),
            .in1(N__1157),
            .in2(N__956),
            .in3(N__808),
            .lcout(signal_out_fsm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1406),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_RNI7RPG_1_LC_14_15_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNI7RPG_1_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNI7RPG_1_LC_14_15_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNI7RPG_1_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__1070),
            .in2(_gnd_net_),
            .in3(N__807),
            .lcout(\fsm_shiftRegs_inst1.un1_current_state4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_RNO_1_2_LC_14_15_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_1_2_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_1_2_LC_14_15_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNO_1_2_LC_14_15_3  (
            .in0(N__1071),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1043),
            .lcout(\fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.en_fin_LC_15_13_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.en_fin_LC_15_13_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.en_fin_LC_15_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fsm_shiftRegs_inst1.en_fin_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__955),
            .lcout(ENdin_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1414),
            .ce(),
            .sr(N__1372));
    defparam \fsm_shiftRegs_inst1.current_state_3_LC_15_14_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_3_LC_15_14_0 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.current_state_3_LC_15_14_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_3_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__993),
            .in2(_gnd_net_),
            .in3(N__962),
            .lcout(\fsm_shiftRegs_inst1.current_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1412),
            .ce(),
            .sr(N__1370));
    defparam \fsm_shiftRegs_inst1.sel_dyn_LC_15_14_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.sel_dyn_LC_15_14_3 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.sel_dyn_LC_15_14_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \fsm_shiftRegs_inst1.sel_dyn_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__951),
            .in2(_gnd_net_),
            .in3(N__1262),
            .lcout(SELDYN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1412),
            .ce(),
            .sr(N__1370));
    defparam \fsm_shiftRegs_inst1.bit_sequence_10_LC_15_15_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_10_LC_15_15_0 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_10_LC_15_15_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_10_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__1302),
            .in2(_gnd_net_),
            .in3(N__1133),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1409),
            .ce(N__1090),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_11_LC_15_15_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_11_LC_15_15_1 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_11_LC_15_15_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_11_LC_15_15_1  (
            .in0(N__1303),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__911),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1409),
            .ce(N__1090),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_13_LC_15_15_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_13_LC_15_15_2 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_13_LC_15_15_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_13_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(N__1305),
            .in2(_gnd_net_),
            .in3(N__1145),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1409),
            .ce(N__1090),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_14_LC_15_15_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_14_LC_15_15_3 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_14_LC_15_15_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_14_LC_15_15_3  (
            .in0(N__1306),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__905),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1409),
            .ce(N__1090),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_8_LC_15_15_4 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_8_LC_15_15_4 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_8_LC_15_15_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_8_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(N__1308),
            .in2(_gnd_net_),
            .in3(N__1121),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1409),
            .ce(N__1090),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_15_LC_15_15_5 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_15_LC_15_15_5 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_15_LC_15_15_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_15_LC_15_15_5  (
            .in0(N__1307),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1163),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1409),
            .ce(N__1090),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_12_LC_15_15_6 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_12_LC_15_15_6 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_12_LC_15_15_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_12_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(N__1304),
            .in2(_gnd_net_),
            .in3(N__1151),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1409),
            .ce(N__1090),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_9_LC_15_15_7 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_9_LC_15_15_7 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_9_LC_15_15_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_9_LC_15_15_7  (
            .in0(N__1309),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1139),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1409),
            .ce(N__1090),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_6_LC_15_16_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_6_LC_15_16_0 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_6_LC_15_16_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_6_LC_15_16_0  (
            .in0(_gnd_net_),
            .in1(N__1313),
            .in2(_gnd_net_),
            .in3(N__1097),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1407),
            .ce(N__1091),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_2_LC_15_16_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_2_LC_15_16_1 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_2_LC_15_16_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_2_LC_15_16_1  (
            .in0(N__1315),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1407),
            .ce(N__1091),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_7_LC_15_16_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_7_LC_15_16_3 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_7_LC_15_16_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_7_LC_15_16_3  (
            .in0(N__1314),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1127),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1407),
            .ce(N__1091),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_3_LC_15_16_4 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_3_LC_15_16_4 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_3_LC_15_16_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_3_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(N__1310),
            .in2(_gnd_net_),
            .in3(N__1115),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1407),
            .ce(N__1091),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_4_LC_15_16_5 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_4_LC_15_16_5 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_4_LC_15_16_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_4_LC_15_16_5  (
            .in0(N__1311),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1109),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1407),
            .ce(N__1091),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_5_LC_15_16_6 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_5_LC_15_16_6 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_5_LC_15_16_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_5_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(N__1312),
            .in2(_gnd_net_),
            .in3(N__1103),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1407),
            .ce(N__1091),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.sel_stat_LC_16_14_6 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.sel_stat_LC_16_14_6 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.sel_stat_LC_16_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fsm_shiftRegs_inst1.sel_stat_LC_16_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1340),
            .lcout(SELSTAT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1415),
            .ce(),
            .sr(N__1373));
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_4_LC_16_15_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_4_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_4_LC_16_15_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNO_0_4_LC_16_15_0  (
            .in0(N__1553),
            .in1(N__1180),
            .in2(N__1580),
            .in3(N__1516),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_4_LC_16_15_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_4_LC_16_15_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.current_state_4_LC_16_15_1 .LUT_INIT=16'b1100111011101110;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_4_LC_16_15_1  (
            .in0(N__1260),
            .in1(N__1339),
            .in2(N__1328),
            .in3(N__1241),
            .lcout(\fsm_shiftRegs_inst1.current_stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1413),
            .ce(),
            .sr(N__1371));
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_0_LC_16_15_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_0_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_0_LC_16_15_2 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNO_0_0_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(N__1552),
            .in2(N__1579),
            .in3(N__1515),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_0_LC_16_15_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_0_LC_16_15_3 .SEQ_MODE=4'b1011;
    defparam \fsm_shiftRegs_inst1.current_state_0_LC_16_15_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_0_LC_16_15_3  (
            .in0(N__1181),
            .in1(N__1261),
            .in2(N__1325),
            .in3(N__1240),
            .lcout(\fsm_shiftRegs_inst1.current_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1413),
            .ce(),
            .sr(N__1371));
    defparam \fsm_shiftRegs_inst1.current_state_RNIVA94_4_LC_16_15_4 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNIVA94_4_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNIVA94_4_LC_16_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNIVA94_4_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1259),
            .lcout(\fsm_shiftRegs_inst1.current_state_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counter2_RNITAO81_7_LC_16_15_5 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter2_RNITAO81_7_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.counter2_RNITAO81_7_LC_16_15_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_RNITAO81_7_LC_16_15_5  (
            .in0(N__1495),
            .in1(N__1531),
            .in2(N__1481),
            .in3(N__1426),
            .lcout(\fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.signal_aux_LC_16_15_7 .C_ON=1'b0;
    defparam \generator_inst1.signal_aux_LC_16_15_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.signal_aux_LC_16_15_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \generator_inst1.signal_aux_LC_16_15_7  (
            .in0(N__1232),
            .in1(N__1226),
            .in2(_gnd_net_),
            .in3(N__1211),
            .lcout(generated_signal_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1413),
            .ce(),
            .sr(N__1371));
    defparam \fsm_shiftRegs_inst1.counter2_0_LC_16_16_0 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_0_LC_16_16_0 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_0_LC_16_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_0_LC_16_16_0  (
            .in0(N__1457),
            .in1(N__1179),
            .in2(_gnd_net_),
            .in3(N__1166),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_0 ),
            .ltout(),
            .carryin(bfn_16_16_0_),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_0 ),
            .clk(N__1410),
            .ce(),
            .sr(N__1367));
    defparam \fsm_shiftRegs_inst1.counter2_1_LC_16_16_1 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_1_LC_16_16_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_1_LC_16_16_1 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_1_LC_16_16_1  (
            .in0(N__1453),
            .in1(_gnd_net_),
            .in2(N__1578),
            .in3(N__1556),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_1 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_0 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_1 ),
            .clk(N__1410),
            .ce(),
            .sr(N__1367));
    defparam \fsm_shiftRegs_inst1.counter2_2_LC_16_16_2 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_2_LC_16_16_2 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_2_LC_16_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_2_LC_16_16_2  (
            .in0(N__1458),
            .in1(N__1551),
            .in2(_gnd_net_),
            .in3(N__1535),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_2 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_1 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_2 ),
            .clk(N__1410),
            .ce(),
            .sr(N__1367));
    defparam \fsm_shiftRegs_inst1.counter2_3_LC_16_16_3 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_3_LC_16_16_3 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_3_LC_16_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_3_LC_16_16_3  (
            .in0(N__1454),
            .in1(N__1532),
            .in2(_gnd_net_),
            .in3(N__1520),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_3 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_2 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_3 ),
            .clk(N__1410),
            .ce(),
            .sr(N__1367));
    defparam \fsm_shiftRegs_inst1.counter2_4_LC_16_16_4 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_4_LC_16_16_4 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_4_LC_16_16_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_4_LC_16_16_4  (
            .in0(N__1459),
            .in1(_gnd_net_),
            .in2(N__1517),
            .in3(N__1499),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_4 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_3 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_4 ),
            .clk(N__1410),
            .ce(),
            .sr(N__1367));
    defparam \fsm_shiftRegs_inst1.counter2_5_LC_16_16_5 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_5_LC_16_16_5 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_5_LC_16_16_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_5_LC_16_16_5  (
            .in0(N__1455),
            .in1(N__1496),
            .in2(_gnd_net_),
            .in3(N__1484),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_5 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_4 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_5 ),
            .clk(N__1410),
            .ce(),
            .sr(N__1367));
    defparam \fsm_shiftRegs_inst1.counter2_6_LC_16_16_6 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_6_LC_16_16_6 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_6_LC_16_16_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_6_LC_16_16_6  (
            .in0(N__1460),
            .in1(N__1477),
            .in2(_gnd_net_),
            .in3(N__1463),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_6 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_5 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_6 ),
            .clk(N__1410),
            .ce(),
            .sr(N__1367));
    defparam \fsm_shiftRegs_inst1.counter2_7_LC_16_16_7 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter2_7_LC_16_16_7 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_7_LC_16_16_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_7_LC_16_16_7  (
            .in0(N__1456),
            .in1(N__1427),
            .in2(_gnd_net_),
            .in3(N__1430),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1410),
            .ce(),
            .sr(N__1367));
endmodule // top
