-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 18 2025 10:14:08

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    generated_signal : out std_logic;
    RST_N : in std_logic;
    ENdin : out std_logic;
    CLK : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__1640\ : std_logic;
signal \N__1639\ : std_logic;
signal \N__1638\ : std_logic;
signal \N__1629\ : std_logic;
signal \N__1628\ : std_logic;
signal \N__1627\ : std_logic;
signal \N__1620\ : std_logic;
signal \N__1619\ : std_logic;
signal \N__1618\ : std_logic;
signal \N__1611\ : std_logic;
signal \N__1610\ : std_logic;
signal \N__1609\ : std_logic;
signal \N__1592\ : std_logic;
signal \N__1589\ : std_logic;
signal \N__1588\ : std_logic;
signal \N__1587\ : std_logic;
signal \N__1584\ : std_logic;
signal \N__1581\ : std_logic;
signal \N__1578\ : std_logic;
signal \N__1571\ : std_logic;
signal \N__1568\ : std_logic;
signal \N__1565\ : std_logic;
signal \N__1564\ : std_logic;
signal \N__1563\ : std_logic;
signal \N__1558\ : std_logic;
signal \N__1555\ : std_logic;
signal \N__1550\ : std_logic;
signal \N__1547\ : std_logic;
signal \N__1546\ : std_logic;
signal \N__1543\ : std_logic;
signal \N__1540\ : std_logic;
signal \N__1535\ : std_logic;
signal \N__1532\ : std_logic;
signal \N__1531\ : std_logic;
signal \N__1530\ : std_logic;
signal \N__1527\ : std_logic;
signal \N__1522\ : std_logic;
signal \N__1519\ : std_logic;
signal \N__1514\ : std_logic;
signal \N__1511\ : std_logic;
signal \N__1510\ : std_logic;
signal \N__1507\ : std_logic;
signal \N__1504\ : std_logic;
signal \N__1499\ : std_logic;
signal \N__1496\ : std_logic;
signal \N__1495\ : std_logic;
signal \N__1492\ : std_logic;
signal \N__1489\ : std_logic;
signal \N__1486\ : std_logic;
signal \N__1481\ : std_logic;
signal \N__1478\ : std_logic;
signal \N__1477\ : std_logic;
signal \N__1476\ : std_logic;
signal \N__1475\ : std_logic;
signal \N__1474\ : std_logic;
signal \N__1473\ : std_logic;
signal \N__1472\ : std_logic;
signal \N__1471\ : std_logic;
signal \N__1462\ : std_logic;
signal \N__1453\ : std_logic;
signal \N__1448\ : std_logic;
signal \N__1445\ : std_logic;
signal \N__1444\ : std_logic;
signal \N__1441\ : std_logic;
signal \N__1438\ : std_logic;
signal \N__1433\ : std_logic;
signal \N__1432\ : std_logic;
signal \N__1431\ : std_logic;
signal \N__1430\ : std_logic;
signal \N__1429\ : std_logic;
signal \N__1428\ : std_logic;
signal \N__1427\ : std_logic;
signal \N__1426\ : std_logic;
signal \N__1425\ : std_logic;
signal \N__1424\ : std_logic;
signal \N__1423\ : std_logic;
signal \N__1422\ : std_logic;
signal \N__1397\ : std_logic;
signal \N__1394\ : std_logic;
signal \N__1391\ : std_logic;
signal \N__1390\ : std_logic;
signal \N__1389\ : std_logic;
signal \N__1388\ : std_logic;
signal \N__1387\ : std_logic;
signal \N__1386\ : std_logic;
signal \N__1385\ : std_logic;
signal \N__1384\ : std_logic;
signal \N__1367\ : std_logic;
signal \N__1364\ : std_logic;
signal \N__1361\ : std_logic;
signal \N__1358\ : std_logic;
signal \N__1355\ : std_logic;
signal \N__1352\ : std_logic;
signal \N__1349\ : std_logic;
signal \N__1346\ : std_logic;
signal \N__1343\ : std_logic;
signal \N__1340\ : std_logic;
signal \N__1337\ : std_logic;
signal \N__1334\ : std_logic;
signal \N__1331\ : std_logic;
signal \N__1328\ : std_logic;
signal \N__1325\ : std_logic;
signal \N__1322\ : std_logic;
signal \N__1319\ : std_logic;
signal \N__1318\ : std_logic;
signal \N__1317\ : std_logic;
signal \N__1316\ : std_logic;
signal \N__1315\ : std_logic;
signal \N__1314\ : std_logic;
signal \N__1313\ : std_logic;
signal \N__1310\ : std_logic;
signal \N__1297\ : std_logic;
signal \N__1296\ : std_logic;
signal \N__1295\ : std_logic;
signal \N__1294\ : std_logic;
signal \N__1293\ : std_logic;
signal \N__1292\ : std_logic;
signal \N__1291\ : std_logic;
signal \N__1290\ : std_logic;
signal \N__1289\ : std_logic;
signal \N__1286\ : std_logic;
signal \N__1283\ : std_logic;
signal \N__1266\ : std_logic;
signal \N__1259\ : std_logic;
signal \N__1256\ : std_logic;
signal \N__1253\ : std_logic;
signal \N__1250\ : std_logic;
signal \N__1247\ : std_logic;
signal \N__1246\ : std_logic;
signal \N__1243\ : std_logic;
signal \N__1240\ : std_logic;
signal \N__1235\ : std_logic;
signal \N__1234\ : std_logic;
signal \N__1233\ : std_logic;
signal \N__1228\ : std_logic;
signal \N__1225\ : std_logic;
signal \N__1220\ : std_logic;
signal \N__1217\ : std_logic;
signal \N__1216\ : std_logic;
signal \N__1211\ : std_logic;
signal \N__1208\ : std_logic;
signal \N__1207\ : std_logic;
signal \N__1206\ : std_logic;
signal \N__1205\ : std_logic;
signal \N__1202\ : std_logic;
signal \N__1199\ : std_logic;
signal \N__1194\ : std_logic;
signal \N__1187\ : std_logic;
signal \N__1186\ : std_logic;
signal \N__1183\ : std_logic;
signal \N__1180\ : std_logic;
signal \N__1175\ : std_logic;
signal \N__1172\ : std_logic;
signal \N__1169\ : std_logic;
signal \N__1166\ : std_logic;
signal \N__1163\ : std_logic;
signal \N__1160\ : std_logic;
signal \N__1157\ : std_logic;
signal \N__1154\ : std_logic;
signal \N__1151\ : std_logic;
signal \N__1148\ : std_logic;
signal \N__1145\ : std_logic;
signal \N__1142\ : std_logic;
signal \N__1139\ : std_logic;
signal \N__1136\ : std_logic;
signal \N__1133\ : std_logic;
signal \N__1130\ : std_logic;
signal \N__1127\ : std_logic;
signal \N__1124\ : std_logic;
signal \N__1121\ : std_logic;
signal \N__1118\ : std_logic;
signal \N__1115\ : std_logic;
signal \N__1112\ : std_logic;
signal \N__1109\ : std_logic;
signal \N__1108\ : std_logic;
signal \N__1107\ : std_logic;
signal \N__1106\ : std_logic;
signal \N__1097\ : std_logic;
signal \N__1094\ : std_logic;
signal \N__1093\ : std_logic;
signal \N__1092\ : std_logic;
signal \N__1091\ : std_logic;
signal \N__1090\ : std_logic;
signal \N__1089\ : std_logic;
signal \N__1086\ : std_logic;
signal \N__1083\ : std_logic;
signal \N__1072\ : std_logic;
signal \N__1067\ : std_logic;
signal \N__1066\ : std_logic;
signal \N__1065\ : std_logic;
signal \N__1064\ : std_logic;
signal \N__1061\ : std_logic;
signal \N__1060\ : std_logic;
signal \N__1049\ : std_logic;
signal \N__1046\ : std_logic;
signal \N__1045\ : std_logic;
signal \N__1044\ : std_logic;
signal \N__1043\ : std_logic;
signal \N__1040\ : std_logic;
signal \N__1039\ : std_logic;
signal \N__1036\ : std_logic;
signal \N__1035\ : std_logic;
signal \N__1034\ : std_logic;
signal \N__1033\ : std_logic;
signal \N__1032\ : std_logic;
signal \N__1029\ : std_logic;
signal \N__1026\ : std_logic;
signal \N__1023\ : std_logic;
signal \N__1010\ : std_logic;
signal \N__1001\ : std_logic;
signal \N__1000\ : std_logic;
signal \N__997\ : std_logic;
signal \N__994\ : std_logic;
signal \N__993\ : std_logic;
signal \N__990\ : std_logic;
signal \N__985\ : std_logic;
signal \N__982\ : std_logic;
signal \N__979\ : std_logic;
signal \N__976\ : std_logic;
signal \N__973\ : std_logic;
signal \N__970\ : std_logic;
signal \N__967\ : std_logic;
signal \N__964\ : std_logic;
signal \N__961\ : std_logic;
signal \N__956\ : std_logic;
signal \N__955\ : std_logic;
signal \N__954\ : std_logic;
signal \N__953\ : std_logic;
signal \N__952\ : std_logic;
signal \N__947\ : std_logic;
signal \N__946\ : std_logic;
signal \N__945\ : std_logic;
signal \N__942\ : std_logic;
signal \N__937\ : std_logic;
signal \N__934\ : std_logic;
signal \N__929\ : std_logic;
signal \N__920\ : std_logic;
signal \N__919\ : std_logic;
signal \N__918\ : std_logic;
signal \N__917\ : std_logic;
signal \N__914\ : std_logic;
signal \N__909\ : std_logic;
signal \N__906\ : std_logic;
signal \N__899\ : std_logic;
signal \N__896\ : std_logic;
signal \N__893\ : std_logic;
signal \N__892\ : std_logic;
signal \N__889\ : std_logic;
signal \N__886\ : std_logic;
signal \N__881\ : std_logic;
signal \N__878\ : std_logic;
signal \N__875\ : std_logic;
signal \N__872\ : std_logic;
signal \N__869\ : std_logic;
signal \N__866\ : std_logic;
signal \N__863\ : std_logic;
signal \N__860\ : std_logic;
signal \N__857\ : std_logic;
signal \N__854\ : std_logic;
signal \N__851\ : std_logic;
signal \N__848\ : std_logic;
signal \N__845\ : std_logic;
signal \N__842\ : std_logic;
signal \N__841\ : std_logic;
signal \N__838\ : std_logic;
signal \N__835\ : std_logic;
signal \N__830\ : std_logic;
signal \N__827\ : std_logic;
signal \N__826\ : std_logic;
signal \N__825\ : std_logic;
signal \N__822\ : std_logic;
signal \N__817\ : std_logic;
signal \N__814\ : std_logic;
signal \N__809\ : std_logic;
signal \N__806\ : std_logic;
signal \N__803\ : std_logic;
signal \N__800\ : std_logic;
signal \N__799\ : std_logic;
signal \N__798\ : std_logic;
signal \N__797\ : std_logic;
signal \N__796\ : std_logic;
signal \N__791\ : std_logic;
signal \N__784\ : std_logic;
signal \N__779\ : std_logic;
signal \N__778\ : std_logic;
signal \N__777\ : std_logic;
signal \N__776\ : std_logic;
signal \N__769\ : std_logic;
signal \N__766\ : std_logic;
signal \N__763\ : std_logic;
signal \N__758\ : std_logic;
signal \N__755\ : std_logic;
signal \N__754\ : std_logic;
signal \N__753\ : std_logic;
signal \N__750\ : std_logic;
signal \N__749\ : std_logic;
signal \N__746\ : std_logic;
signal \N__743\ : std_logic;
signal \N__742\ : std_logic;
signal \N__737\ : std_logic;
signal \N__730\ : std_logic;
signal \N__725\ : std_logic;
signal \N__722\ : std_logic;
signal \N__719\ : std_logic;
signal \N__716\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \RST_N_c_i\ : std_logic;
signal \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.counterZ0Z_0\ : std_logic;
signal \fsm_shiftRegs_inst1.counterZ0Z_1\ : std_logic;
signal \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.counterZ0Z_3\ : std_logic;
signal \ENdin_c\ : std_logic;
signal enable_din : std_logic;
signal \fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.N_123_1\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.counterDYNZ0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.counterDYNZ0Z_2\ : std_logic;
signal \fsm_shiftRegs_inst1.counterDYNZ0Z_0\ : std_logic;
signal \fsm_shiftRegs_inst1.counterDYNZ0Z_1\ : std_logic;
signal \fsm_shiftRegs_inst1.current_stateZ0Z_2\ : std_logic;
signal \RST_N_c\ : std_logic;
signal \fsm_shiftRegs_inst1.current_stateZ0Z_1\ : std_logic;
signal \fsm_shiftRegs_inst1.counterZ0Z_2\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2\ : std_logic;
signal \fsm_shiftRegs_inst1.current_stateZ0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0\ : std_logic;
signal \fsm_shiftRegs_inst1.current_stateZ0Z_4\ : std_logic;
signal signal_out_fsm : std_logic;
signal \SELSTAT\ : std_logic;
signal \SELDYN\ : std_logic;
signal generated_signal_c : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_2\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_6\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_4\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_5\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_15\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_11\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_12\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_10\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_13\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_14\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_9\ : std_logic;
signal \fsm_shiftRegs_inst1.current_stateZ0Z_0\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_7\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_8\ : std_logic;
signal \fsm_shiftRegs_inst1.un1_current_state4_0\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_0\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_1\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_0\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_2\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_1\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_2\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_4\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_3\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_5\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_4\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_6\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_5\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_i_4\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_6\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_7\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \CLK_c_g\ : std_logic;
signal \RST_N_c_i_g\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \RST_N_wire\ : std_logic;
signal generated_signal_wire : std_logic;
signal \ENdin_wire\ : std_logic;

begin
    \CLK_wire\ <= CLK;
    \RST_N_wire\ <= RST_N;
    generated_signal <= generated_signal_wire;
    ENdin <= \ENdin_wire\;

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__1638\,
            GLOBALBUFFEROUTPUT => \CLK_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1640\,
            DIN => \N__1639\,
            DOUT => \N__1638\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1640\,
            PADOUT => \N__1639\,
            PADIN => \N__1638\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RST_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1629\,
            DIN => \N__1628\,
            DOUT => \N__1627\,
            PACKAGEPIN => \RST_N_wire\
        );

    \RST_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1629\,
            PADOUT => \N__1628\,
            PADIN => \N__1627\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RST_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \generated_signal_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1620\,
            DIN => \N__1619\,
            DOUT => \N__1618\,
            PACKAGEPIN => generated_signal_wire
        );

    \generated_signal_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1620\,
            PADOUT => \N__1619\,
            PADIN => \N__1618\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1163\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ENdin_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1611\,
            DIN => \N__1610\,
            DOUT => \N__1609\,
            PACKAGEPIN => \ENdin_wire\
        );

    \ENdin_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1611\,
            PADOUT => \N__1610\,
            PADIN => \N__1609\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__875\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__355\ : InMux
    port map (
            O => \N__1592\,
            I => \N__1589\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__1589\,
            I => \N__1584\
        );

    \I__353\ : InMux
    port map (
            O => \N__1588\,
            I => \N__1581\
        );

    \I__352\ : InMux
    port map (
            O => \N__1587\,
            I => \N__1578\
        );

    \I__351\ : Odrv4
    port map (
            O => \N__1584\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_1\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__1581\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_1\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__1578\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_1\
        );

    \I__348\ : InMux
    port map (
            O => \N__1571\,
            I => \fsm_shiftRegs_inst1.counter2_cry_0\
        );

    \I__347\ : CascadeMux
    port map (
            O => \N__1568\,
            I => \N__1565\
        );

    \I__346\ : InMux
    port map (
            O => \N__1565\,
            I => \N__1558\
        );

    \I__345\ : InMux
    port map (
            O => \N__1564\,
            I => \N__1558\
        );

    \I__344\ : InMux
    port map (
            O => \N__1563\,
            I => \N__1555\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__1558\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_2\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__1555\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_2\
        );

    \I__341\ : InMux
    port map (
            O => \N__1550\,
            I => \fsm_shiftRegs_inst1.counter2_cry_1\
        );

    \I__340\ : InMux
    port map (
            O => \N__1547\,
            I => \N__1543\
        );

    \I__339\ : InMux
    port map (
            O => \N__1546\,
            I => \N__1540\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__1543\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_3\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__1540\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_3\
        );

    \I__336\ : InMux
    port map (
            O => \N__1535\,
            I => \fsm_shiftRegs_inst1.counter2_cry_2\
        );

    \I__335\ : CascadeMux
    port map (
            O => \N__1532\,
            I => \N__1527\
        );

    \I__334\ : InMux
    port map (
            O => \N__1531\,
            I => \N__1522\
        );

    \I__333\ : InMux
    port map (
            O => \N__1530\,
            I => \N__1522\
        );

    \I__332\ : InMux
    port map (
            O => \N__1527\,
            I => \N__1519\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__1522\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_4\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__1519\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_4\
        );

    \I__329\ : InMux
    port map (
            O => \N__1514\,
            I => \fsm_shiftRegs_inst1.counter2_cry_3\
        );

    \I__328\ : InMux
    port map (
            O => \N__1511\,
            I => \N__1507\
        );

    \I__327\ : InMux
    port map (
            O => \N__1510\,
            I => \N__1504\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__1507\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_5\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__1504\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_5\
        );

    \I__324\ : InMux
    port map (
            O => \N__1499\,
            I => \fsm_shiftRegs_inst1.counter2_cry_4\
        );

    \I__323\ : CascadeMux
    port map (
            O => \N__1496\,
            I => \N__1492\
        );

    \I__322\ : InMux
    port map (
            O => \N__1495\,
            I => \N__1489\
        );

    \I__321\ : InMux
    port map (
            O => \N__1492\,
            I => \N__1486\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__1489\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_6\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__1486\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_6\
        );

    \I__318\ : InMux
    port map (
            O => \N__1481\,
            I => \fsm_shiftRegs_inst1.counter2_cry_5\
        );

    \I__317\ : InMux
    port map (
            O => \N__1478\,
            I => \N__1462\
        );

    \I__316\ : InMux
    port map (
            O => \N__1477\,
            I => \N__1462\
        );

    \I__315\ : InMux
    port map (
            O => \N__1476\,
            I => \N__1462\
        );

    \I__314\ : InMux
    port map (
            O => \N__1475\,
            I => \N__1462\
        );

    \I__313\ : InMux
    port map (
            O => \N__1474\,
            I => \N__1453\
        );

    \I__312\ : InMux
    port map (
            O => \N__1473\,
            I => \N__1453\
        );

    \I__311\ : InMux
    port map (
            O => \N__1472\,
            I => \N__1453\
        );

    \I__310\ : InMux
    port map (
            O => \N__1471\,
            I => \N__1453\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__1462\,
            I => \fsm_shiftRegs_inst1.current_state_i_4\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__1453\,
            I => \fsm_shiftRegs_inst1.current_state_i_4\
        );

    \I__307\ : InMux
    port map (
            O => \N__1448\,
            I => \fsm_shiftRegs_inst1.counter2_cry_6\
        );

    \I__306\ : InMux
    port map (
            O => \N__1445\,
            I => \N__1441\
        );

    \I__305\ : InMux
    port map (
            O => \N__1444\,
            I => \N__1438\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__1441\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_7\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__1438\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_7\
        );

    \I__302\ : ClkMux
    port map (
            O => \N__1433\,
            I => \N__1397\
        );

    \I__301\ : ClkMux
    port map (
            O => \N__1432\,
            I => \N__1397\
        );

    \I__300\ : ClkMux
    port map (
            O => \N__1431\,
            I => \N__1397\
        );

    \I__299\ : ClkMux
    port map (
            O => \N__1430\,
            I => \N__1397\
        );

    \I__298\ : ClkMux
    port map (
            O => \N__1429\,
            I => \N__1397\
        );

    \I__297\ : ClkMux
    port map (
            O => \N__1428\,
            I => \N__1397\
        );

    \I__296\ : ClkMux
    port map (
            O => \N__1427\,
            I => \N__1397\
        );

    \I__295\ : ClkMux
    port map (
            O => \N__1426\,
            I => \N__1397\
        );

    \I__294\ : ClkMux
    port map (
            O => \N__1425\,
            I => \N__1397\
        );

    \I__293\ : ClkMux
    port map (
            O => \N__1424\,
            I => \N__1397\
        );

    \I__292\ : ClkMux
    port map (
            O => \N__1423\,
            I => \N__1397\
        );

    \I__291\ : ClkMux
    port map (
            O => \N__1422\,
            I => \N__1397\
        );

    \I__290\ : GlobalMux
    port map (
            O => \N__1397\,
            I => \N__1394\
        );

    \I__289\ : gio2CtrlBuf
    port map (
            O => \N__1394\,
            I => \CLK_c_g\
        );

    \I__288\ : SRMux
    port map (
            O => \N__1391\,
            I => \N__1367\
        );

    \I__287\ : SRMux
    port map (
            O => \N__1390\,
            I => \N__1367\
        );

    \I__286\ : SRMux
    port map (
            O => \N__1389\,
            I => \N__1367\
        );

    \I__285\ : SRMux
    port map (
            O => \N__1388\,
            I => \N__1367\
        );

    \I__284\ : SRMux
    port map (
            O => \N__1387\,
            I => \N__1367\
        );

    \I__283\ : SRMux
    port map (
            O => \N__1386\,
            I => \N__1367\
        );

    \I__282\ : SRMux
    port map (
            O => \N__1385\,
            I => \N__1367\
        );

    \I__281\ : SRMux
    port map (
            O => \N__1384\,
            I => \N__1367\
        );

    \I__280\ : GlobalMux
    port map (
            O => \N__1367\,
            I => \N__1364\
        );

    \I__279\ : gio2CtrlBuf
    port map (
            O => \N__1364\,
            I => \RST_N_c_i_g\
        );

    \I__278\ : InMux
    port map (
            O => \N__1361\,
            I => \N__1358\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__1358\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_15\
        );

    \I__276\ : InMux
    port map (
            O => \N__1355\,
            I => \N__1352\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__1352\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_11\
        );

    \I__274\ : InMux
    port map (
            O => \N__1349\,
            I => \N__1346\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__1346\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_12\
        );

    \I__272\ : InMux
    port map (
            O => \N__1343\,
            I => \N__1340\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__1340\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_10\
        );

    \I__270\ : InMux
    port map (
            O => \N__1337\,
            I => \N__1334\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__1334\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_13\
        );

    \I__268\ : InMux
    port map (
            O => \N__1331\,
            I => \N__1328\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__1328\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_14\
        );

    \I__266\ : InMux
    port map (
            O => \N__1325\,
            I => \N__1322\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__1322\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_9\
        );

    \I__264\ : CascadeMux
    port map (
            O => \N__1319\,
            I => \N__1310\
        );

    \I__263\ : InMux
    port map (
            O => \N__1318\,
            I => \N__1297\
        );

    \I__262\ : InMux
    port map (
            O => \N__1317\,
            I => \N__1297\
        );

    \I__261\ : InMux
    port map (
            O => \N__1316\,
            I => \N__1297\
        );

    \I__260\ : InMux
    port map (
            O => \N__1315\,
            I => \N__1297\
        );

    \I__259\ : InMux
    port map (
            O => \N__1314\,
            I => \N__1297\
        );

    \I__258\ : InMux
    port map (
            O => \N__1313\,
            I => \N__1297\
        );

    \I__257\ : InMux
    port map (
            O => \N__1310\,
            I => \N__1286\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__1297\,
            I => \N__1283\
        );

    \I__255\ : InMux
    port map (
            O => \N__1296\,
            I => \N__1266\
        );

    \I__254\ : InMux
    port map (
            O => \N__1295\,
            I => \N__1266\
        );

    \I__253\ : InMux
    port map (
            O => \N__1294\,
            I => \N__1266\
        );

    \I__252\ : InMux
    port map (
            O => \N__1293\,
            I => \N__1266\
        );

    \I__251\ : InMux
    port map (
            O => \N__1292\,
            I => \N__1266\
        );

    \I__250\ : InMux
    port map (
            O => \N__1291\,
            I => \N__1266\
        );

    \I__249\ : InMux
    port map (
            O => \N__1290\,
            I => \N__1266\
        );

    \I__248\ : InMux
    port map (
            O => \N__1289\,
            I => \N__1266\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__1286\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_0\
        );

    \I__246\ : Odrv4
    port map (
            O => \N__1283\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_0\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__1266\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_0\
        );

    \I__244\ : InMux
    port map (
            O => \N__1259\,
            I => \N__1256\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__1256\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_7\
        );

    \I__242\ : InMux
    port map (
            O => \N__1253\,
            I => \N__1250\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__1250\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_8\
        );

    \I__240\ : CEMux
    port map (
            O => \N__1247\,
            I => \N__1243\
        );

    \I__239\ : CEMux
    port map (
            O => \N__1246\,
            I => \N__1240\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__1243\,
            I => \fsm_shiftRegs_inst1.un1_current_state4_0\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__1240\,
            I => \fsm_shiftRegs_inst1.un1_current_state4_0\
        );

    \I__236\ : InMux
    port map (
            O => \N__1235\,
            I => \N__1228\
        );

    \I__235\ : InMux
    port map (
            O => \N__1234\,
            I => \N__1228\
        );

    \I__234\ : InMux
    port map (
            O => \N__1233\,
            I => \N__1225\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__1228\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_0\
        );

    \I__232\ : LocalMux
    port map (
            O => \N__1225\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_0\
        );

    \I__231\ : InMux
    port map (
            O => \N__1220\,
            I => \bfn_14_15_0_\
        );

    \I__230\ : InMux
    port map (
            O => \N__1217\,
            I => \N__1211\
        );

    \I__229\ : InMux
    port map (
            O => \N__1216\,
            I => \N__1211\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__1211\,
            I => \fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0\
        );

    \I__227\ : InMux
    port map (
            O => \N__1208\,
            I => \N__1202\
        );

    \I__226\ : InMux
    port map (
            O => \N__1207\,
            I => \N__1199\
        );

    \I__225\ : InMux
    port map (
            O => \N__1206\,
            I => \N__1194\
        );

    \I__224\ : InMux
    port map (
            O => \N__1205\,
            I => \N__1194\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__1202\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_4\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__1199\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_4\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__1194\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_4\
        );

    \I__220\ : InMux
    port map (
            O => \N__1187\,
            I => \N__1183\
        );

    \I__219\ : InMux
    port map (
            O => \N__1186\,
            I => \N__1180\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__1183\,
            I => signal_out_fsm
        );

    \I__217\ : LocalMux
    port map (
            O => \N__1180\,
            I => signal_out_fsm
        );

    \I__216\ : InMux
    port map (
            O => \N__1175\,
            I => \N__1172\
        );

    \I__215\ : LocalMux
    port map (
            O => \N__1172\,
            I => \SELSTAT\
        );

    \I__214\ : InMux
    port map (
            O => \N__1169\,
            I => \N__1166\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__1166\,
            I => \SELDYN\
        );

    \I__212\ : IoInMux
    port map (
            O => \N__1163\,
            I => \N__1160\
        );

    \I__211\ : LocalMux
    port map (
            O => \N__1160\,
            I => \N__1157\
        );

    \I__210\ : Span4Mux_s1_v
    port map (
            O => \N__1157\,
            I => \N__1154\
        );

    \I__209\ : Span4Mux_v
    port map (
            O => \N__1154\,
            I => \N__1151\
        );

    \I__208\ : Sp12to4
    port map (
            O => \N__1151\,
            I => \N__1148\
        );

    \I__207\ : Span12Mux_s10_h
    port map (
            O => \N__1148\,
            I => \N__1145\
        );

    \I__206\ : Span12Mux_v
    port map (
            O => \N__1145\,
            I => \N__1142\
        );

    \I__205\ : Odrv12
    port map (
            O => \N__1142\,
            I => generated_signal_c
        );

    \I__204\ : InMux
    port map (
            O => \N__1139\,
            I => \N__1136\
        );

    \I__203\ : LocalMux
    port map (
            O => \N__1136\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_2\
        );

    \I__202\ : InMux
    port map (
            O => \N__1133\,
            I => \N__1130\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__1130\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_3\
        );

    \I__200\ : InMux
    port map (
            O => \N__1127\,
            I => \N__1124\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__1124\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_6\
        );

    \I__198\ : InMux
    port map (
            O => \N__1121\,
            I => \N__1118\
        );

    \I__197\ : LocalMux
    port map (
            O => \N__1118\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_4\
        );

    \I__196\ : InMux
    port map (
            O => \N__1115\,
            I => \N__1112\
        );

    \I__195\ : LocalMux
    port map (
            O => \N__1112\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_5\
        );

    \I__194\ : InMux
    port map (
            O => \N__1109\,
            I => \N__1097\
        );

    \I__193\ : InMux
    port map (
            O => \N__1108\,
            I => \N__1097\
        );

    \I__192\ : InMux
    port map (
            O => \N__1107\,
            I => \N__1097\
        );

    \I__191\ : InMux
    port map (
            O => \N__1106\,
            I => \N__1097\
        );

    \I__190\ : LocalMux
    port map (
            O => \N__1097\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_2\
        );

    \I__189\ : CascadeMux
    port map (
            O => \N__1094\,
            I => \N__1086\
        );

    \I__188\ : InMux
    port map (
            O => \N__1093\,
            I => \N__1083\
        );

    \I__187\ : InMux
    port map (
            O => \N__1092\,
            I => \N__1072\
        );

    \I__186\ : InMux
    port map (
            O => \N__1091\,
            I => \N__1072\
        );

    \I__185\ : InMux
    port map (
            O => \N__1090\,
            I => \N__1072\
        );

    \I__184\ : InMux
    port map (
            O => \N__1089\,
            I => \N__1072\
        );

    \I__183\ : InMux
    port map (
            O => \N__1086\,
            I => \N__1072\
        );

    \I__182\ : LocalMux
    port map (
            O => \N__1083\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_0\
        );

    \I__181\ : LocalMux
    port map (
            O => \N__1072\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_0\
        );

    \I__180\ : CascadeMux
    port map (
            O => \N__1067\,
            I => \N__1061\
        );

    \I__179\ : InMux
    port map (
            O => \N__1066\,
            I => \N__1049\
        );

    \I__178\ : InMux
    port map (
            O => \N__1065\,
            I => \N__1049\
        );

    \I__177\ : InMux
    port map (
            O => \N__1064\,
            I => \N__1049\
        );

    \I__176\ : InMux
    port map (
            O => \N__1061\,
            I => \N__1049\
        );

    \I__175\ : InMux
    port map (
            O => \N__1060\,
            I => \N__1049\
        );

    \I__174\ : LocalMux
    port map (
            O => \N__1049\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_1\
        );

    \I__173\ : InMux
    port map (
            O => \N__1046\,
            I => \N__1040\
        );

    \I__172\ : CascadeMux
    port map (
            O => \N__1045\,
            I => \N__1036\
        );

    \I__171\ : InMux
    port map (
            O => \N__1044\,
            I => \N__1029\
        );

    \I__170\ : InMux
    port map (
            O => \N__1043\,
            I => \N__1026\
        );

    \I__169\ : LocalMux
    port map (
            O => \N__1040\,
            I => \N__1023\
        );

    \I__168\ : InMux
    port map (
            O => \N__1039\,
            I => \N__1010\
        );

    \I__167\ : InMux
    port map (
            O => \N__1036\,
            I => \N__1010\
        );

    \I__166\ : InMux
    port map (
            O => \N__1035\,
            I => \N__1010\
        );

    \I__165\ : InMux
    port map (
            O => \N__1034\,
            I => \N__1010\
        );

    \I__164\ : InMux
    port map (
            O => \N__1033\,
            I => \N__1010\
        );

    \I__163\ : InMux
    port map (
            O => \N__1032\,
            I => \N__1010\
        );

    \I__162\ : LocalMux
    port map (
            O => \N__1029\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_2\
        );

    \I__161\ : LocalMux
    port map (
            O => \N__1026\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_2\
        );

    \I__160\ : Odrv4
    port map (
            O => \N__1023\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_2\
        );

    \I__159\ : LocalMux
    port map (
            O => \N__1010\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_2\
        );

    \I__158\ : InMux
    port map (
            O => \N__1001\,
            I => \N__997\
        );

    \I__157\ : CascadeMux
    port map (
            O => \N__1000\,
            I => \N__994\
        );

    \I__156\ : LocalMux
    port map (
            O => \N__997\,
            I => \N__990\
        );

    \I__155\ : InMux
    port map (
            O => \N__994\,
            I => \N__985\
        );

    \I__154\ : InMux
    port map (
            O => \N__993\,
            I => \N__985\
        );

    \I__153\ : Sp12to4
    port map (
            O => \N__990\,
            I => \N__982\
        );

    \I__152\ : LocalMux
    port map (
            O => \N__985\,
            I => \N__979\
        );

    \I__151\ : Span12Mux_v
    port map (
            O => \N__982\,
            I => \N__976\
        );

    \I__150\ : Sp12to4
    port map (
            O => \N__979\,
            I => \N__973\
        );

    \I__149\ : Span12Mux_h
    port map (
            O => \N__976\,
            I => \N__970\
        );

    \I__148\ : Span12Mux_v
    port map (
            O => \N__973\,
            I => \N__967\
        );

    \I__147\ : Span12Mux_h
    port map (
            O => \N__970\,
            I => \N__964\
        );

    \I__146\ : Span12Mux_h
    port map (
            O => \N__967\,
            I => \N__961\
        );

    \I__145\ : Odrv12
    port map (
            O => \N__964\,
            I => \RST_N_c\
        );

    \I__144\ : Odrv12
    port map (
            O => \N__961\,
            I => \RST_N_c\
        );

    \I__143\ : InMux
    port map (
            O => \N__956\,
            I => \N__947\
        );

    \I__142\ : InMux
    port map (
            O => \N__955\,
            I => \N__947\
        );

    \I__141\ : InMux
    port map (
            O => \N__954\,
            I => \N__942\
        );

    \I__140\ : InMux
    port map (
            O => \N__953\,
            I => \N__937\
        );

    \I__139\ : InMux
    port map (
            O => \N__952\,
            I => \N__937\
        );

    \I__138\ : LocalMux
    port map (
            O => \N__947\,
            I => \N__934\
        );

    \I__137\ : InMux
    port map (
            O => \N__946\,
            I => \N__929\
        );

    \I__136\ : InMux
    port map (
            O => \N__945\,
            I => \N__929\
        );

    \I__135\ : LocalMux
    port map (
            O => \N__942\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_1\
        );

    \I__134\ : LocalMux
    port map (
            O => \N__937\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_1\
        );

    \I__133\ : Odrv4
    port map (
            O => \N__934\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_1\
        );

    \I__132\ : LocalMux
    port map (
            O => \N__929\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_1\
        );

    \I__131\ : InMux
    port map (
            O => \N__920\,
            I => \N__914\
        );

    \I__130\ : InMux
    port map (
            O => \N__919\,
            I => \N__909\
        );

    \I__129\ : InMux
    port map (
            O => \N__918\,
            I => \N__909\
        );

    \I__128\ : InMux
    port map (
            O => \N__917\,
            I => \N__906\
        );

    \I__127\ : LocalMux
    port map (
            O => \N__914\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_2\
        );

    \I__126\ : LocalMux
    port map (
            O => \N__909\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_2\
        );

    \I__125\ : LocalMux
    port map (
            O => \N__906\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_2\
        );

    \I__124\ : InMux
    port map (
            O => \N__899\,
            I => \N__896\
        );

    \I__123\ : LocalMux
    port map (
            O => \N__896\,
            I => \fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2\
        );

    \I__122\ : InMux
    port map (
            O => \N__893\,
            I => \N__889\
        );

    \I__121\ : InMux
    port map (
            O => \N__892\,
            I => \N__886\
        );

    \I__120\ : LocalMux
    port map (
            O => \N__889\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_3\
        );

    \I__119\ : LocalMux
    port map (
            O => \N__886\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_3\
        );

    \I__118\ : CascadeMux
    port map (
            O => \N__881\,
            I => \fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_\
        );

    \I__117\ : CascadeMux
    port map (
            O => \N__878\,
            I => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_\
        );

    \I__116\ : IoInMux
    port map (
            O => \N__875\,
            I => \N__872\
        );

    \I__115\ : LocalMux
    port map (
            O => \N__872\,
            I => \N__869\
        );

    \I__114\ : IoSpan4Mux
    port map (
            O => \N__869\,
            I => \N__866\
        );

    \I__113\ : Sp12to4
    port map (
            O => \N__866\,
            I => \N__863\
        );

    \I__112\ : Span12Mux_s7_h
    port map (
            O => \N__863\,
            I => \N__860\
        );

    \I__111\ : Span12Mux_h
    port map (
            O => \N__860\,
            I => \N__857\
        );

    \I__110\ : Odrv12
    port map (
            O => \N__857\,
            I => \ENdin_c\
        );

    \I__109\ : InMux
    port map (
            O => \N__854\,
            I => \N__851\
        );

    \I__108\ : LocalMux
    port map (
            O => \N__851\,
            I => enable_din
        );

    \I__107\ : CascadeMux
    port map (
            O => \N__848\,
            I => \fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_\
        );

    \I__106\ : InMux
    port map (
            O => \N__845\,
            I => \N__842\
        );

    \I__105\ : LocalMux
    port map (
            O => \N__842\,
            I => \N__838\
        );

    \I__104\ : InMux
    port map (
            O => \N__841\,
            I => \N__835\
        );

    \I__103\ : Odrv4
    port map (
            O => \N__838\,
            I => \fsm_shiftRegs_inst1.N_123_1\
        );

    \I__102\ : LocalMux
    port map (
            O => \N__835\,
            I => \fsm_shiftRegs_inst1.N_123_1\
        );

    \I__101\ : CascadeMux
    port map (
            O => \N__830\,
            I => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_\
        );

    \I__100\ : CascadeMux
    port map (
            O => \N__827\,
            I => \N__822\
        );

    \I__99\ : InMux
    port map (
            O => \N__826\,
            I => \N__817\
        );

    \I__98\ : InMux
    port map (
            O => \N__825\,
            I => \N__817\
        );

    \I__97\ : InMux
    port map (
            O => \N__822\,
            I => \N__814\
        );

    \I__96\ : LocalMux
    port map (
            O => \N__817\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_3\
        );

    \I__95\ : LocalMux
    port map (
            O => \N__814\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_3\
        );

    \I__94\ : InMux
    port map (
            O => \N__809\,
            I => \N__806\
        );

    \I__93\ : LocalMux
    port map (
            O => \N__806\,
            I => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3\
        );

    \I__92\ : CascadeMux
    port map (
            O => \N__803\,
            I => \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_\
        );

    \I__91\ : InMux
    port map (
            O => \N__800\,
            I => \N__791\
        );

    \I__90\ : InMux
    port map (
            O => \N__799\,
            I => \N__791\
        );

    \I__89\ : InMux
    port map (
            O => \N__798\,
            I => \N__784\
        );

    \I__88\ : InMux
    port map (
            O => \N__797\,
            I => \N__784\
        );

    \I__87\ : InMux
    port map (
            O => \N__796\,
            I => \N__784\
        );

    \I__86\ : LocalMux
    port map (
            O => \N__791\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_0\
        );

    \I__85\ : LocalMux
    port map (
            O => \N__784\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_0\
        );

    \I__84\ : InMux
    port map (
            O => \N__779\,
            I => \N__769\
        );

    \I__83\ : InMux
    port map (
            O => \N__778\,
            I => \N__769\
        );

    \I__82\ : InMux
    port map (
            O => \N__777\,
            I => \N__769\
        );

    \I__81\ : InMux
    port map (
            O => \N__776\,
            I => \N__766\
        );

    \I__80\ : LocalMux
    port map (
            O => \N__769\,
            I => \N__763\
        );

    \I__79\ : LocalMux
    port map (
            O => \N__766\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_1\
        );

    \I__78\ : Odrv4
    port map (
            O => \N__763\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_1\
        );

    \I__77\ : CascadeMux
    port map (
            O => \N__758\,
            I => \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3_cascade_\
        );

    \I__76\ : CascadeMux
    port map (
            O => \N__755\,
            I => \N__750\
        );

    \I__75\ : CascadeMux
    port map (
            O => \N__754\,
            I => \N__746\
        );

    \I__74\ : CascadeMux
    port map (
            O => \N__753\,
            I => \N__743\
        );

    \I__73\ : InMux
    port map (
            O => \N__750\,
            I => \N__737\
        );

    \I__72\ : InMux
    port map (
            O => \N__749\,
            I => \N__737\
        );

    \I__71\ : InMux
    port map (
            O => \N__746\,
            I => \N__730\
        );

    \I__70\ : InMux
    port map (
            O => \N__743\,
            I => \N__730\
        );

    \I__69\ : InMux
    port map (
            O => \N__742\,
            I => \N__730\
        );

    \I__68\ : LocalMux
    port map (
            O => \N__737\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_3\
        );

    \I__67\ : LocalMux
    port map (
            O => \N__730\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_3\
        );

    \I__66\ : IoInMux
    port map (
            O => \N__725\,
            I => \N__722\
        );

    \I__65\ : LocalMux
    port map (
            O => \N__722\,
            I => \N__719\
        );

    \I__64\ : Span4Mux_s3_h
    port map (
            O => \N__719\,
            I => \N__716\
        );

    \I__63\ : Odrv4
    port map (
            O => \N__716\,
            I => \RST_N_c_i\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_15_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \RST_N_ibuf_RNIBJGC_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__725\,
            GLOBALBUFFEROUTPUT => \RST_N_c_i_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \RST_N_ibuf_RNIBJGC_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1001\,
            lcout => \RST_N_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counter_0_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__955\,
            in1 => \N__749\,
            in2 => \_gnd_net_\,
            in3 => \N__800\,
            lcout => \fsm_shiftRegs_inst1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1423\,
            ce => 'H',
            sr => \N__1385\
        );

    \fsm_shiftRegs_inst1.counter_1_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100010000001000"
        )
    port map (
            in0 => \N__799\,
            in1 => \N__956\,
            in2 => \N__755\,
            in3 => \N__776\,
            lcout => \fsm_shiftRegs_inst1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1423\,
            ce => 'H',
            sr => \N__1385\
        );

    \fsm_shiftRegs_inst1.counter_RNO_0_2_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100001000"
        )
    port map (
            in0 => \N__797\,
            in1 => \N__778\,
            in2 => \N__753\,
            in3 => \N__918\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counter_2_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__952\,
            in1 => \_gnd_net_\,
            in2 => \N__803\,
            in3 => \_gnd_net_\,
            lcout => \fsm_shiftRegs_inst1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1426\,
            ce => 'H',
            sr => \N__1388\
        );

    \fsm_shiftRegs_inst1.counter_RNIC589_1_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__777\,
            in1 => \N__796\,
            in2 => \_gnd_net_\,
            in3 => \N__742\,
            lcout => \fsm_shiftRegs_inst1.N_123_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counter_RNO_0_3_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__798\,
            in1 => \N__779\,
            in2 => \N__754\,
            in3 => \N__919\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counter_3_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__953\,
            in1 => \_gnd_net_\,
            in2 => \N__758\,
            in3 => \_gnd_net_\,
            lcout => \fsm_shiftRegs_inst1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1426\,
            ce => 'H',
            sr => \N__1388\
        );

    \fsm_shiftRegs_inst1.current_state_1_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011111010"
        )
    port map (
            in0 => \N__954\,
            in1 => \N__920\,
            in2 => \N__1319\,
            in3 => \N__841\,
            lcout => \fsm_shiftRegs_inst1.current_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1424\,
            ce => 'H',
            sr => \N__1386\
        );

    \fsm_shiftRegs_inst1.current_state_3_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1093\,
            in2 => \_gnd_net_\,
            in3 => \N__809\,
            lcout => \fsm_shiftRegs_inst1.current_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1424\,
            ce => 'H',
            sr => \N__1386\
        );

    \fsm_shiftRegs_inst1.sel_stat_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__893\,
            lcout => \SELSTAT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1422\,
            ce => 'H',
            sr => \N__1384\
        );

    \fsm_shiftRegs_inst1.sel_dyn_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1046\,
            in2 => \_gnd_net_\,
            in3 => \N__1208\,
            lcout => \SELDYN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1422\,
            ce => 'H',
            sr => \N__1384\
        );

    \enableDin_aux_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__854\,
            lcout => \ENdin_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.en_fin_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1044\,
            lcout => enable_din,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1431\,
            ce => 'H',
            sr => \N__1391\
        );

    \fsm_shiftRegs_inst1.counterDYN_RNO_0_3_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__825\,
            in1 => \N__1089\,
            in2 => \N__1067\,
            in3 => \N__1108\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counterDYN_3_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__848\,
            in3 => \N__1039\,
            lcout => \fsm_shiftRegs_inst1.counterDYNZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1429\,
            ce => 'H',
            sr => \N__1390\
        );

    \fsm_shiftRegs_inst1.counterDYN_0_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__1033\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1091\,
            lcout => \fsm_shiftRegs_inst1.counterDYNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1429\,
            ce => 'H',
            sr => \N__1390\
        );

    \fsm_shiftRegs_inst1.current_state_RNO_0_2_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__1107\,
            in1 => \N__1064\,
            in2 => \N__1094\,
            in3 => \N__826\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_2_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__1034\,
            in1 => \N__845\,
            in2 => \N__830\,
            in3 => \N__899\,
            lcout => \fsm_shiftRegs_inst1.current_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1429\,
            ce => 'H',
            sr => \N__1390\
        );

    \fsm_shiftRegs_inst1.current_state_RNO_0_3_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1106\,
            in1 => \N__1060\,
            in2 => \N__827\,
            in3 => \N__1032\,
            lcout => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counterDYN_2_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000010000000"
        )
    port map (
            in0 => \N__1065\,
            in1 => \N__1092\,
            in2 => \N__1045\,
            in3 => \N__1109\,
            lcout => \fsm_shiftRegs_inst1.counterDYNZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1429\,
            ce => 'H',
            sr => \N__1390\
        );

    \fsm_shiftRegs_inst1.counterDYN_1_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__1090\,
            in1 => \N__1035\,
            in2 => \_gnd_net_\,
            in3 => \N__1066\,
            lcout => \fsm_shiftRegs_inst1.counterDYNZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1429\,
            ce => 'H',
            sr => \N__1390\
        );

    \fsm_shiftRegs_inst1.signal_out_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__1187\,
            in1 => \N__1361\,
            in2 => \N__1000\,
            in3 => \N__1043\,
            lcout => signal_out_fsm,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_RNI7RPG_1_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__993\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__945\,
            lcout => \fsm_shiftRegs_inst1.un1_current_state4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_RNO_1_2_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__946\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__917\,
            lcout => \fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_RNO_0_4_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__1592\,
            in1 => \N__1234\,
            in2 => \N__1568\,
            in3 => \N__1531\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_4_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111011101110"
        )
    port map (
            in0 => \N__1207\,
            in1 => \N__892\,
            in2 => \N__881\,
            in3 => \N__1217\,
            lcout => \fsm_shiftRegs_inst1.current_stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1425\,
            ce => 'H',
            sr => \N__1387\
        );

    \fsm_shiftRegs_inst1.current_state_RNO_0_0_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__1564\,
            in1 => \N__1588\,
            in2 => \_gnd_net_\,
            in3 => \N__1530\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_0_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__1235\,
            in1 => \N__1206\,
            in2 => \N__878\,
            in3 => \N__1216\,
            lcout => \fsm_shiftRegs_inst1.current_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1425\,
            ce => 'H',
            sr => \N__1387\
        );

    \fsm_shiftRegs_inst1.counter2_RNITAO81_7_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1510\,
            in1 => \N__1546\,
            in2 => \N__1496\,
            in3 => \N__1444\,
            lcout => \fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_RNIVA94_4_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1205\,
            lcout => \fsm_shiftRegs_inst1.current_state_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.signal_aux_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__1186\,
            in1 => \N__1175\,
            in2 => \_gnd_net_\,
            in3 => \N__1169\,
            lcout => generated_signal_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1425\,
            ce => 'H',
            sr => \N__1387\
        );

    \fsm_shiftRegs_inst1.bit_sequence_3_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1313\,
            in2 => \_gnd_net_\,
            in3 => \N__1139\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1432\,
            ce => \N__1247\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_2_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__1318\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1432\,
            ce => \N__1247\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_4_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1314\,
            in2 => \_gnd_net_\,
            in3 => \N__1133\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1432\,
            ce => \N__1247\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_6_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__1316\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1115\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1432\,
            ce => \N__1247\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_7_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1317\,
            in2 => \_gnd_net_\,
            in3 => \N__1127\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1432\,
            ce => \N__1247\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_5_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__1315\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1121\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1432\,
            ce => \N__1247\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_15_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1294\,
            in2 => \_gnd_net_\,
            in3 => \N__1331\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1430\,
            ce => \N__1246\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_11_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__1290\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1343\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1430\,
            ce => \N__1246\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_12_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1291\,
            in2 => \_gnd_net_\,
            in3 => \N__1355\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1430\,
            ce => \N__1246\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_13_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__1292\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1349\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1430\,
            ce => \N__1246\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_10_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1289\,
            in2 => \_gnd_net_\,
            in3 => \N__1325\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1430\,
            ce => \N__1246\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_14_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__1293\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1337\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1430\,
            ce => \N__1246\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_9_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1296\,
            in2 => \_gnd_net_\,
            in3 => \N__1253\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1430\,
            ce => \N__1246\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_8_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__1295\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1259\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1430\,
            ce => \N__1246\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counter2_0_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1475\,
            in1 => \N__1233\,
            in2 => \_gnd_net_\,
            in3 => \N__1220\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_0\,
            clk => \N__1428\,
            ce => 'H',
            sr => \N__1389\
        );

    \fsm_shiftRegs_inst1.counter2_1_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1471\,
            in1 => \N__1587\,
            in2 => \_gnd_net_\,
            in3 => \N__1571\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_1\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_0\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_1\,
            clk => \N__1428\,
            ce => 'H',
            sr => \N__1389\
        );

    \fsm_shiftRegs_inst1.counter2_2_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1476\,
            in1 => \N__1563\,
            in2 => \_gnd_net_\,
            in3 => \N__1550\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_2\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_1\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_2\,
            clk => \N__1428\,
            ce => 'H',
            sr => \N__1389\
        );

    \fsm_shiftRegs_inst1.counter2_3_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1472\,
            in1 => \N__1547\,
            in2 => \_gnd_net_\,
            in3 => \N__1535\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_3\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_2\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_3\,
            clk => \N__1428\,
            ce => 'H',
            sr => \N__1389\
        );

    \fsm_shiftRegs_inst1.counter2_4_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__1477\,
            in1 => \_gnd_net_\,
            in2 => \N__1532\,
            in3 => \N__1514\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_4\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_3\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_4\,
            clk => \N__1428\,
            ce => 'H',
            sr => \N__1389\
        );

    \fsm_shiftRegs_inst1.counter2_5_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1473\,
            in1 => \N__1511\,
            in2 => \_gnd_net_\,
            in3 => \N__1499\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_5\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_4\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_5\,
            clk => \N__1428\,
            ce => 'H',
            sr => \N__1389\
        );

    \fsm_shiftRegs_inst1.counter2_6_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1478\,
            in1 => \N__1495\,
            in2 => \_gnd_net_\,
            in3 => \N__1481\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_6\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_5\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_6\,
            clk => \N__1428\,
            ce => 'H',
            sr => \N__1389\
        );

    \fsm_shiftRegs_inst1.counter2_7_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1474\,
            in1 => \N__1445\,
            in2 => \_gnd_net_\,
            in3 => \N__1448\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1428\,
            ce => 'H',
            sr => \N__1389\
        );
end \INTERFACE\;
