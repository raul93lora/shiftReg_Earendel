// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 18 2025 08:30:48

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    generated_signal,
    RST_N,
    ENFIN,
    CLK);

    output generated_signal;
    input RST_N;
    output ENFIN;
    input CLK;

    wire N__1656;
    wire N__1655;
    wire N__1654;
    wire N__1645;
    wire N__1644;
    wire N__1643;
    wire N__1636;
    wire N__1635;
    wire N__1634;
    wire N__1627;
    wire N__1626;
    wire N__1625;
    wire N__1608;
    wire N__1605;
    wire N__1602;
    wire N__1601;
    wire N__1600;
    wire N__1595;
    wire N__1592;
    wire N__1587;
    wire N__1584;
    wire N__1583;
    wire N__1580;
    wire N__1577;
    wire N__1572;
    wire N__1569;
    wire N__1568;
    wire N__1567;
    wire N__1564;
    wire N__1559;
    wire N__1556;
    wire N__1551;
    wire N__1548;
    wire N__1547;
    wire N__1544;
    wire N__1541;
    wire N__1538;
    wire N__1533;
    wire N__1530;
    wire N__1527;
    wire N__1526;
    wire N__1523;
    wire N__1520;
    wire N__1515;
    wire N__1512;
    wire N__1509;
    wire N__1508;
    wire N__1505;
    wire N__1502;
    wire N__1497;
    wire N__1496;
    wire N__1495;
    wire N__1494;
    wire N__1493;
    wire N__1492;
    wire N__1491;
    wire N__1490;
    wire N__1489;
    wire N__1488;
    wire N__1487;
    wire N__1464;
    wire N__1461;
    wire N__1458;
    wire N__1457;
    wire N__1456;
    wire N__1455;
    wire N__1454;
    wire N__1453;
    wire N__1452;
    wire N__1437;
    wire N__1434;
    wire N__1431;
    wire N__1430;
    wire N__1429;
    wire N__1428;
    wire N__1425;
    wire N__1422;
    wire N__1421;
    wire N__1418;
    wire N__1415;
    wire N__1412;
    wire N__1409;
    wire N__1406;
    wire N__1395;
    wire N__1394;
    wire N__1393;
    wire N__1392;
    wire N__1391;
    wire N__1390;
    wire N__1389;
    wire N__1388;
    wire N__1379;
    wire N__1370;
    wire N__1365;
    wire N__1364;
    wire N__1361;
    wire N__1358;
    wire N__1355;
    wire N__1350;
    wire N__1347;
    wire N__1344;
    wire N__1343;
    wire N__1338;
    wire N__1335;
    wire N__1334;
    wire N__1333;
    wire N__1332;
    wire N__1331;
    wire N__1330;
    wire N__1329;
    wire N__1328;
    wire N__1327;
    wire N__1326;
    wire N__1323;
    wire N__1320;
    wire N__1317;
    wire N__1314;
    wire N__1305;
    wire N__1300;
    wire N__1287;
    wire N__1286;
    wire N__1283;
    wire N__1280;
    wire N__1277;
    wire N__1274;
    wire N__1269;
    wire N__1268;
    wire N__1267;
    wire N__1264;
    wire N__1263;
    wire N__1260;
    wire N__1257;
    wire N__1254;
    wire N__1251;
    wire N__1248;
    wire N__1245;
    wire N__1240;
    wire N__1235;
    wire N__1232;
    wire N__1229;
    wire N__1224;
    wire N__1223;
    wire N__1222;
    wire N__1221;
    wire N__1220;
    wire N__1219;
    wire N__1218;
    wire N__1217;
    wire N__1216;
    wire N__1215;
    wire N__1214;
    wire N__1213;
    wire N__1212;
    wire N__1211;
    wire N__1210;
    wire N__1207;
    wire N__1206;
    wire N__1205;
    wire N__1202;
    wire N__1187;
    wire N__1174;
    wire N__1171;
    wire N__1166;
    wire N__1155;
    wire N__1154;
    wire N__1151;
    wire N__1148;
    wire N__1143;
    wire N__1140;
    wire N__1137;
    wire N__1134;
    wire N__1133;
    wire N__1132;
    wire N__1127;
    wire N__1124;
    wire N__1119;
    wire N__1116;
    wire N__1113;
    wire N__1112;
    wire N__1111;
    wire N__1108;
    wire N__1105;
    wire N__1102;
    wire N__1095;
    wire N__1092;
    wire N__1089;
    wire N__1086;
    wire N__1083;
    wire N__1080;
    wire N__1077;
    wire N__1074;
    wire N__1071;
    wire N__1068;
    wire N__1065;
    wire N__1062;
    wire N__1059;
    wire N__1056;
    wire N__1053;
    wire N__1050;
    wire N__1047;
    wire N__1046;
    wire N__1045;
    wire N__1044;
    wire N__1041;
    wire N__1040;
    wire N__1039;
    wire N__1036;
    wire N__1027;
    wire N__1024;
    wire N__1017;
    wire N__1014;
    wire N__1011;
    wire N__1010;
    wire N__1009;
    wire N__1008;
    wire N__1005;
    wire N__1002;
    wire N__1001;
    wire N__996;
    wire N__989;
    wire N__984;
    wire N__983;
    wire N__982;
    wire N__981;
    wire N__980;
    wire N__977;
    wire N__976;
    wire N__973;
    wire N__970;
    wire N__961;
    wire N__954;
    wire N__953;
    wire N__952;
    wire N__951;
    wire N__950;
    wire N__947;
    wire N__944;
    wire N__937;
    wire N__934;
    wire N__927;
    wire N__924;
    wire N__923;
    wire N__922;
    wire N__921;
    wire N__918;
    wire N__911;
    wire N__906;
    wire N__903;
    wire N__900;
    wire N__897;
    wire N__894;
    wire N__891;
    wire N__888;
    wire N__885;
    wire N__882;
    wire N__879;
    wire N__876;
    wire N__873;
    wire N__870;
    wire N__867;
    wire N__864;
    wire N__861;
    wire N__858;
    wire N__857;
    wire N__856;
    wire N__855;
    wire N__854;
    wire N__851;
    wire N__842;
    wire N__837;
    wire N__836;
    wire N__835;
    wire N__834;
    wire N__831;
    wire N__824;
    wire N__819;
    wire N__816;
    wire N__815;
    wire N__814;
    wire N__813;
    wire N__810;
    wire N__803;
    wire N__798;
    wire N__795;
    wire N__792;
    wire N__789;
    wire N__786;
    wire N__783;
    wire N__780;
    wire N__779;
    wire N__776;
    wire N__775;
    wire N__768;
    wire N__765;
    wire N__762;
    wire N__759;
    wire N__758;
    wire N__755;
    wire N__752;
    wire N__747;
    wire N__744;
    wire N__741;
    wire N__738;
    wire N__735;
    wire N__732;
    wire N__729;
    wire N__726;
    wire N__723;
    wire N__720;
    wire N__717;
    wire VCCG0;
    wire GNDG0;
    wire signal_out_fsm;
    wire SELSTAT;
    wire SELDYN;
    wire generated_signal_c;
    wire RST_N_c_i;
    wire \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_ ;
    wire \fsm_shiftRegs_inst1.N_125_1_cascade_ ;
    wire \fsm_shiftRegs_inst1.counterZ0Z_0 ;
    wire \fsm_shiftRegs_inst1.counterZ0Z_1 ;
    wire \fsm_shiftRegs_inst1.counterZ0Z_2 ;
    wire \fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_ ;
    wire \fsm_shiftRegs_inst1.N_125_1 ;
    wire \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_ ;
    wire \fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2 ;
    wire \fsm_shiftRegs_inst1.counterDYNZ0Z_3 ;
    wire \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3 ;
    wire \fsm_shiftRegs_inst1.counterDYNZ0Z_2 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_15 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_14 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_13 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_12 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_11 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_10 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_5 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_6 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_3 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_4 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_7 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_8 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_9 ;
    wire ENFIN_c;
    wire \fsm_shiftRegs_inst1.current_stateZ0Z_1 ;
    wire \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3 ;
    wire \fsm_shiftRegs_inst1.counterZ0Z_3 ;
    wire \fsm_shiftRegs_inst1.counterDYNZ0Z_0 ;
    wire \fsm_shiftRegs_inst1.counterDYNZ0Z_1 ;
    wire \fsm_shiftRegs_inst1.current_stateZ0Z_3 ;
    wire \fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_ ;
    wire \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_ ;
    wire \fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0 ;
    wire \fsm_shiftRegs_inst1.current_stateZ0Z_2 ;
    wire \fsm_shiftRegs_inst1.un1_current_state4_0 ;
    wire RST_N_c;
    wire \fsm_shiftRegs_inst1.current_stateZ0Z_0 ;
    wire \fsm_shiftRegs_inst1.bit_sequenceZ0Z_2 ;
    wire \fsm_shiftRegs_inst1.N_122_i ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_0 ;
    wire bfn_4_11_0_;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_1 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_0 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_2 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_1 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_3 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_2 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_4 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_3 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_5 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_4 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_6 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_5 ;
    wire \fsm_shiftRegs_inst1.counter2_cry_6 ;
    wire \fsm_shiftRegs_inst1.counter2Z0Z_7 ;
    wire CLK_c_g;
    wire RST_N_c_i_g;
    wire \fsm_shiftRegs_inst1.current_stateZ0Z_4 ;
    wire \fsm_shiftRegs_inst1.current_state_i_4 ;
    wire _gnd_net_;

    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__1654),
            .GLOBALBUFFEROUTPUT(CLK_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__1656),
            .DIN(N__1655),
            .DOUT(N__1654),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__1656),
            .PADOUT(N__1655),
            .PADIN(N__1654),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RST_N_ibuf_iopad (
            .OE(N__1645),
            .DIN(N__1644),
            .DOUT(N__1643),
            .PACKAGEPIN(RST_N));
    defparam RST_N_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RST_N_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RST_N_ibuf_preio (
            .PADOEN(N__1645),
            .PADOUT(N__1644),
            .PADIN(N__1643),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RST_N_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ENFIN_obuf_iopad (
            .OE(N__1636),
            .DIN(N__1635),
            .DOUT(N__1634),
            .PACKAGEPIN(ENFIN));
    defparam ENFIN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ENFIN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ENFIN_obuf_preio (
            .PADOEN(N__1636),
            .PADOUT(N__1635),
            .PADIN(N__1634),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1059),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD generated_signal_obuf_iopad (
            .OE(N__1627),
            .DIN(N__1626),
            .DOUT(N__1625),
            .PACKAGEPIN(generated_signal));
    defparam generated_signal_obuf_preio.NEG_TRIGGER=1'b0;
    defparam generated_signal_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO generated_signal_obuf_preio (
            .PADOEN(N__1627),
            .PADOUT(N__1626),
            .PADIN(N__1625),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__735),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__360 (
            .O(N__1608),
            .I(\fsm_shiftRegs_inst1.counter2_cry_0 ));
    CascadeMux I__359 (
            .O(N__1605),
            .I(N__1602));
    InMux I__358 (
            .O(N__1602),
            .I(N__1595));
    InMux I__357 (
            .O(N__1601),
            .I(N__1595));
    InMux I__356 (
            .O(N__1600),
            .I(N__1592));
    LocalMux I__355 (
            .O(N__1595),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_2 ));
    LocalMux I__354 (
            .O(N__1592),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_2 ));
    InMux I__353 (
            .O(N__1587),
            .I(\fsm_shiftRegs_inst1.counter2_cry_1 ));
    InMux I__352 (
            .O(N__1584),
            .I(N__1580));
    InMux I__351 (
            .O(N__1583),
            .I(N__1577));
    LocalMux I__350 (
            .O(N__1580),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_3 ));
    LocalMux I__349 (
            .O(N__1577),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_3 ));
    InMux I__348 (
            .O(N__1572),
            .I(\fsm_shiftRegs_inst1.counter2_cry_2 ));
    CascadeMux I__347 (
            .O(N__1569),
            .I(N__1564));
    InMux I__346 (
            .O(N__1568),
            .I(N__1559));
    InMux I__345 (
            .O(N__1567),
            .I(N__1559));
    InMux I__344 (
            .O(N__1564),
            .I(N__1556));
    LocalMux I__343 (
            .O(N__1559),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_4 ));
    LocalMux I__342 (
            .O(N__1556),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_4 ));
    InMux I__341 (
            .O(N__1551),
            .I(\fsm_shiftRegs_inst1.counter2_cry_3 ));
    CascadeMux I__340 (
            .O(N__1548),
            .I(N__1544));
    InMux I__339 (
            .O(N__1547),
            .I(N__1541));
    InMux I__338 (
            .O(N__1544),
            .I(N__1538));
    LocalMux I__337 (
            .O(N__1541),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_5 ));
    LocalMux I__336 (
            .O(N__1538),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_5 ));
    InMux I__335 (
            .O(N__1533),
            .I(\fsm_shiftRegs_inst1.counter2_cry_4 ));
    CascadeMux I__334 (
            .O(N__1530),
            .I(N__1527));
    InMux I__333 (
            .O(N__1527),
            .I(N__1523));
    InMux I__332 (
            .O(N__1526),
            .I(N__1520));
    LocalMux I__331 (
            .O(N__1523),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_6 ));
    LocalMux I__330 (
            .O(N__1520),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_6 ));
    InMux I__329 (
            .O(N__1515),
            .I(\fsm_shiftRegs_inst1.counter2_cry_5 ));
    InMux I__328 (
            .O(N__1512),
            .I(\fsm_shiftRegs_inst1.counter2_cry_6 ));
    InMux I__327 (
            .O(N__1509),
            .I(N__1505));
    InMux I__326 (
            .O(N__1508),
            .I(N__1502));
    LocalMux I__325 (
            .O(N__1505),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_7 ));
    LocalMux I__324 (
            .O(N__1502),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_7 ));
    ClkMux I__323 (
            .O(N__1497),
            .I(N__1464));
    ClkMux I__322 (
            .O(N__1496),
            .I(N__1464));
    ClkMux I__321 (
            .O(N__1495),
            .I(N__1464));
    ClkMux I__320 (
            .O(N__1494),
            .I(N__1464));
    ClkMux I__319 (
            .O(N__1493),
            .I(N__1464));
    ClkMux I__318 (
            .O(N__1492),
            .I(N__1464));
    ClkMux I__317 (
            .O(N__1491),
            .I(N__1464));
    ClkMux I__316 (
            .O(N__1490),
            .I(N__1464));
    ClkMux I__315 (
            .O(N__1489),
            .I(N__1464));
    ClkMux I__314 (
            .O(N__1488),
            .I(N__1464));
    ClkMux I__313 (
            .O(N__1487),
            .I(N__1464));
    GlobalMux I__312 (
            .O(N__1464),
            .I(N__1461));
    gio2CtrlBuf I__311 (
            .O(N__1461),
            .I(CLK_c_g));
    SRMux I__310 (
            .O(N__1458),
            .I(N__1437));
    SRMux I__309 (
            .O(N__1457),
            .I(N__1437));
    SRMux I__308 (
            .O(N__1456),
            .I(N__1437));
    SRMux I__307 (
            .O(N__1455),
            .I(N__1437));
    SRMux I__306 (
            .O(N__1454),
            .I(N__1437));
    SRMux I__305 (
            .O(N__1453),
            .I(N__1437));
    SRMux I__304 (
            .O(N__1452),
            .I(N__1437));
    GlobalMux I__303 (
            .O(N__1437),
            .I(N__1434));
    gio2CtrlBuf I__302 (
            .O(N__1434),
            .I(RST_N_c_i_g));
    InMux I__301 (
            .O(N__1431),
            .I(N__1425));
    InMux I__300 (
            .O(N__1430),
            .I(N__1422));
    InMux I__299 (
            .O(N__1429),
            .I(N__1418));
    InMux I__298 (
            .O(N__1428),
            .I(N__1415));
    LocalMux I__297 (
            .O(N__1425),
            .I(N__1412));
    LocalMux I__296 (
            .O(N__1422),
            .I(N__1409));
    InMux I__295 (
            .O(N__1421),
            .I(N__1406));
    LocalMux I__294 (
            .O(N__1418),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_4 ));
    LocalMux I__293 (
            .O(N__1415),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_4 ));
    Odrv4 I__292 (
            .O(N__1412),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_4 ));
    Odrv4 I__291 (
            .O(N__1409),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_4 ));
    LocalMux I__290 (
            .O(N__1406),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_4 ));
    InMux I__289 (
            .O(N__1395),
            .I(N__1379));
    InMux I__288 (
            .O(N__1394),
            .I(N__1379));
    InMux I__287 (
            .O(N__1393),
            .I(N__1379));
    InMux I__286 (
            .O(N__1392),
            .I(N__1379));
    InMux I__285 (
            .O(N__1391),
            .I(N__1370));
    InMux I__284 (
            .O(N__1390),
            .I(N__1370));
    InMux I__283 (
            .O(N__1389),
            .I(N__1370));
    InMux I__282 (
            .O(N__1388),
            .I(N__1370));
    LocalMux I__281 (
            .O(N__1379),
            .I(\fsm_shiftRegs_inst1.current_state_i_4 ));
    LocalMux I__280 (
            .O(N__1370),
            .I(\fsm_shiftRegs_inst1.current_state_i_4 ));
    InMux I__279 (
            .O(N__1365),
            .I(N__1361));
    InMux I__278 (
            .O(N__1364),
            .I(N__1358));
    LocalMux I__277 (
            .O(N__1361),
            .I(N__1355));
    LocalMux I__276 (
            .O(N__1358),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_3 ));
    Odrv12 I__275 (
            .O(N__1355),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_3 ));
    CascadeMux I__274 (
            .O(N__1350),
            .I(\fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_ ));
    CascadeMux I__273 (
            .O(N__1347),
            .I(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_ ));
    InMux I__272 (
            .O(N__1344),
            .I(N__1338));
    InMux I__271 (
            .O(N__1343),
            .I(N__1338));
    LocalMux I__270 (
            .O(N__1338),
            .I(\fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0 ));
    InMux I__269 (
            .O(N__1335),
            .I(N__1323));
    InMux I__268 (
            .O(N__1334),
            .I(N__1320));
    InMux I__267 (
            .O(N__1333),
            .I(N__1317));
    InMux I__266 (
            .O(N__1332),
            .I(N__1314));
    InMux I__265 (
            .O(N__1331),
            .I(N__1305));
    InMux I__264 (
            .O(N__1330),
            .I(N__1305));
    InMux I__263 (
            .O(N__1329),
            .I(N__1305));
    InMux I__262 (
            .O(N__1328),
            .I(N__1305));
    InMux I__261 (
            .O(N__1327),
            .I(N__1300));
    InMux I__260 (
            .O(N__1326),
            .I(N__1300));
    LocalMux I__259 (
            .O(N__1323),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ));
    LocalMux I__258 (
            .O(N__1320),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ));
    LocalMux I__257 (
            .O(N__1317),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ));
    LocalMux I__256 (
            .O(N__1314),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ));
    LocalMux I__255 (
            .O(N__1305),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ));
    LocalMux I__254 (
            .O(N__1300),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ));
    CEMux I__253 (
            .O(N__1287),
            .I(N__1283));
    CEMux I__252 (
            .O(N__1286),
            .I(N__1280));
    LocalMux I__251 (
            .O(N__1283),
            .I(N__1277));
    LocalMux I__250 (
            .O(N__1280),
            .I(N__1274));
    Odrv4 I__249 (
            .O(N__1277),
            .I(\fsm_shiftRegs_inst1.un1_current_state4_0 ));
    Odrv4 I__248 (
            .O(N__1274),
            .I(\fsm_shiftRegs_inst1.un1_current_state4_0 ));
    InMux I__247 (
            .O(N__1269),
            .I(N__1264));
    InMux I__246 (
            .O(N__1268),
            .I(N__1260));
    CascadeMux I__245 (
            .O(N__1267),
            .I(N__1257));
    LocalMux I__244 (
            .O(N__1264),
            .I(N__1254));
    InMux I__243 (
            .O(N__1263),
            .I(N__1251));
    LocalMux I__242 (
            .O(N__1260),
            .I(N__1248));
    InMux I__241 (
            .O(N__1257),
            .I(N__1245));
    Span4Mux_v I__240 (
            .O(N__1254),
            .I(N__1240));
    LocalMux I__239 (
            .O(N__1251),
            .I(N__1240));
    Span4Mux_v I__238 (
            .O(N__1248),
            .I(N__1235));
    LocalMux I__237 (
            .O(N__1245),
            .I(N__1235));
    Span4Mux_v I__236 (
            .O(N__1240),
            .I(N__1232));
    Span4Mux_v I__235 (
            .O(N__1235),
            .I(N__1229));
    Odrv4 I__234 (
            .O(N__1232),
            .I(RST_N_c));
    Odrv4 I__233 (
            .O(N__1229),
            .I(RST_N_c));
    InMux I__232 (
            .O(N__1224),
            .I(N__1207));
    InMux I__231 (
            .O(N__1223),
            .I(N__1202));
    InMux I__230 (
            .O(N__1222),
            .I(N__1187));
    InMux I__229 (
            .O(N__1221),
            .I(N__1187));
    InMux I__228 (
            .O(N__1220),
            .I(N__1187));
    InMux I__227 (
            .O(N__1219),
            .I(N__1187));
    InMux I__226 (
            .O(N__1218),
            .I(N__1187));
    InMux I__225 (
            .O(N__1217),
            .I(N__1187));
    InMux I__224 (
            .O(N__1216),
            .I(N__1187));
    InMux I__223 (
            .O(N__1215),
            .I(N__1174));
    InMux I__222 (
            .O(N__1214),
            .I(N__1174));
    InMux I__221 (
            .O(N__1213),
            .I(N__1174));
    InMux I__220 (
            .O(N__1212),
            .I(N__1174));
    InMux I__219 (
            .O(N__1211),
            .I(N__1174));
    InMux I__218 (
            .O(N__1210),
            .I(N__1174));
    LocalMux I__217 (
            .O(N__1207),
            .I(N__1171));
    InMux I__216 (
            .O(N__1206),
            .I(N__1166));
    InMux I__215 (
            .O(N__1205),
            .I(N__1166));
    LocalMux I__214 (
            .O(N__1202),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_0 ));
    LocalMux I__213 (
            .O(N__1187),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_0 ));
    LocalMux I__212 (
            .O(N__1174),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_0 ));
    Odrv4 I__211 (
            .O(N__1171),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_0 ));
    LocalMux I__210 (
            .O(N__1166),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_0 ));
    InMux I__209 (
            .O(N__1155),
            .I(N__1151));
    InMux I__208 (
            .O(N__1154),
            .I(N__1148));
    LocalMux I__207 (
            .O(N__1151),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_2 ));
    LocalMux I__206 (
            .O(N__1148),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_2 ));
    CEMux I__205 (
            .O(N__1143),
            .I(N__1140));
    LocalMux I__204 (
            .O(N__1140),
            .I(N__1137));
    Odrv12 I__203 (
            .O(N__1137),
            .I(\fsm_shiftRegs_inst1.N_122_i ));
    InMux I__202 (
            .O(N__1134),
            .I(N__1127));
    InMux I__201 (
            .O(N__1133),
            .I(N__1127));
    InMux I__200 (
            .O(N__1132),
            .I(N__1124));
    LocalMux I__199 (
            .O(N__1127),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_0 ));
    LocalMux I__198 (
            .O(N__1124),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_0 ));
    InMux I__197 (
            .O(N__1119),
            .I(bfn_4_11_0_));
    InMux I__196 (
            .O(N__1116),
            .I(N__1113));
    LocalMux I__195 (
            .O(N__1113),
            .I(N__1108));
    InMux I__194 (
            .O(N__1112),
            .I(N__1105));
    InMux I__193 (
            .O(N__1111),
            .I(N__1102));
    Odrv4 I__192 (
            .O(N__1108),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_1 ));
    LocalMux I__191 (
            .O(N__1105),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_1 ));
    LocalMux I__190 (
            .O(N__1102),
            .I(\fsm_shiftRegs_inst1.counter2Z0Z_1 ));
    InMux I__189 (
            .O(N__1095),
            .I(N__1092));
    LocalMux I__188 (
            .O(N__1092),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_6 ));
    InMux I__187 (
            .O(N__1089),
            .I(N__1086));
    LocalMux I__186 (
            .O(N__1086),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_3 ));
    InMux I__185 (
            .O(N__1083),
            .I(N__1080));
    LocalMux I__184 (
            .O(N__1080),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_4 ));
    InMux I__183 (
            .O(N__1077),
            .I(N__1074));
    LocalMux I__182 (
            .O(N__1074),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_7 ));
    InMux I__181 (
            .O(N__1071),
            .I(N__1068));
    LocalMux I__180 (
            .O(N__1068),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_8 ));
    InMux I__179 (
            .O(N__1065),
            .I(N__1062));
    LocalMux I__178 (
            .O(N__1062),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_9 ));
    IoInMux I__177 (
            .O(N__1059),
            .I(N__1056));
    LocalMux I__176 (
            .O(N__1056),
            .I(N__1053));
    Span4Mux_s1_h I__175 (
            .O(N__1053),
            .I(N__1050));
    Odrv4 I__174 (
            .O(N__1050),
            .I(ENFIN_c));
    CascadeMux I__173 (
            .O(N__1047),
            .I(N__1041));
    InMux I__172 (
            .O(N__1046),
            .I(N__1036));
    InMux I__171 (
            .O(N__1045),
            .I(N__1027));
    InMux I__170 (
            .O(N__1044),
            .I(N__1027));
    InMux I__169 (
            .O(N__1041),
            .I(N__1027));
    InMux I__168 (
            .O(N__1040),
            .I(N__1027));
    InMux I__167 (
            .O(N__1039),
            .I(N__1024));
    LocalMux I__166 (
            .O(N__1036),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_1 ));
    LocalMux I__165 (
            .O(N__1027),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_1 ));
    LocalMux I__164 (
            .O(N__1024),
            .I(\fsm_shiftRegs_inst1.current_stateZ0Z_1 ));
    InMux I__163 (
            .O(N__1017),
            .I(N__1014));
    LocalMux I__162 (
            .O(N__1014),
            .I(\fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3 ));
    CascadeMux I__161 (
            .O(N__1011),
            .I(N__1005));
    CascadeMux I__160 (
            .O(N__1010),
            .I(N__1002));
    InMux I__159 (
            .O(N__1009),
            .I(N__996));
    InMux I__158 (
            .O(N__1008),
            .I(N__996));
    InMux I__157 (
            .O(N__1005),
            .I(N__989));
    InMux I__156 (
            .O(N__1002),
            .I(N__989));
    InMux I__155 (
            .O(N__1001),
            .I(N__989));
    LocalMux I__154 (
            .O(N__996),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_3 ));
    LocalMux I__153 (
            .O(N__989),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_3 ));
    CascadeMux I__152 (
            .O(N__984),
            .I(N__977));
    InMux I__151 (
            .O(N__983),
            .I(N__973));
    InMux I__150 (
            .O(N__982),
            .I(N__970));
    InMux I__149 (
            .O(N__981),
            .I(N__961));
    InMux I__148 (
            .O(N__980),
            .I(N__961));
    InMux I__147 (
            .O(N__977),
            .I(N__961));
    InMux I__146 (
            .O(N__976),
            .I(N__961));
    LocalMux I__145 (
            .O(N__973),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_0 ));
    LocalMux I__144 (
            .O(N__970),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_0 ));
    LocalMux I__143 (
            .O(N__961),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_0 ));
    CascadeMux I__142 (
            .O(N__954),
            .I(N__947));
    InMux I__141 (
            .O(N__953),
            .I(N__944));
    InMux I__140 (
            .O(N__952),
            .I(N__937));
    InMux I__139 (
            .O(N__951),
            .I(N__937));
    InMux I__138 (
            .O(N__950),
            .I(N__937));
    InMux I__137 (
            .O(N__947),
            .I(N__934));
    LocalMux I__136 (
            .O(N__944),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_1 ));
    LocalMux I__135 (
            .O(N__937),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_1 ));
    LocalMux I__134 (
            .O(N__934),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_1 ));
    CascadeMux I__133 (
            .O(N__927),
            .I(N__924));
    InMux I__132 (
            .O(N__924),
            .I(N__918));
    InMux I__131 (
            .O(N__923),
            .I(N__911));
    InMux I__130 (
            .O(N__922),
            .I(N__911));
    InMux I__129 (
            .O(N__921),
            .I(N__911));
    LocalMux I__128 (
            .O(N__918),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_2 ));
    LocalMux I__127 (
            .O(N__911),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_2 ));
    InMux I__126 (
            .O(N__906),
            .I(N__903));
    LocalMux I__125 (
            .O(N__903),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_15 ));
    InMux I__124 (
            .O(N__900),
            .I(N__897));
    LocalMux I__123 (
            .O(N__897),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_14 ));
    InMux I__122 (
            .O(N__894),
            .I(N__891));
    LocalMux I__121 (
            .O(N__891),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_13 ));
    InMux I__120 (
            .O(N__888),
            .I(N__885));
    LocalMux I__119 (
            .O(N__885),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_12 ));
    InMux I__118 (
            .O(N__882),
            .I(N__879));
    LocalMux I__117 (
            .O(N__879),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_11 ));
    InMux I__116 (
            .O(N__876),
            .I(N__873));
    LocalMux I__115 (
            .O(N__873),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_10 ));
    InMux I__114 (
            .O(N__870),
            .I(N__867));
    LocalMux I__113 (
            .O(N__867),
            .I(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_5 ));
    CascadeMux I__112 (
            .O(N__864),
            .I(\fsm_shiftRegs_inst1.N_125_1_cascade_ ));
    CascadeMux I__111 (
            .O(N__861),
            .I(N__858));
    InMux I__110 (
            .O(N__858),
            .I(N__851));
    InMux I__109 (
            .O(N__857),
            .I(N__842));
    InMux I__108 (
            .O(N__856),
            .I(N__842));
    InMux I__107 (
            .O(N__855),
            .I(N__842));
    InMux I__106 (
            .O(N__854),
            .I(N__842));
    LocalMux I__105 (
            .O(N__851),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_0 ));
    LocalMux I__104 (
            .O(N__842),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_0 ));
    InMux I__103 (
            .O(N__837),
            .I(N__831));
    InMux I__102 (
            .O(N__836),
            .I(N__824));
    InMux I__101 (
            .O(N__835),
            .I(N__824));
    InMux I__100 (
            .O(N__834),
            .I(N__824));
    LocalMux I__99 (
            .O(N__831),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_1 ));
    LocalMux I__98 (
            .O(N__824),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_1 ));
    CascadeMux I__97 (
            .O(N__819),
            .I(N__816));
    InMux I__96 (
            .O(N__816),
            .I(N__810));
    InMux I__95 (
            .O(N__815),
            .I(N__803));
    InMux I__94 (
            .O(N__814),
            .I(N__803));
    InMux I__93 (
            .O(N__813),
            .I(N__803));
    LocalMux I__92 (
            .O(N__810),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_2 ));
    LocalMux I__91 (
            .O(N__803),
            .I(\fsm_shiftRegs_inst1.counterZ0Z_2 ));
    CascadeMux I__90 (
            .O(N__798),
            .I(\fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_ ));
    InMux I__89 (
            .O(N__795),
            .I(N__792));
    LocalMux I__88 (
            .O(N__792),
            .I(\fsm_shiftRegs_inst1.N_125_1 ));
    CascadeMux I__87 (
            .O(N__789),
            .I(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_ ));
    InMux I__86 (
            .O(N__786),
            .I(N__783));
    LocalMux I__85 (
            .O(N__783),
            .I(\fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2 ));
    CascadeMux I__84 (
            .O(N__780),
            .I(N__776));
    InMux I__83 (
            .O(N__779),
            .I(N__768));
    InMux I__82 (
            .O(N__776),
            .I(N__768));
    InMux I__81 (
            .O(N__775),
            .I(N__768));
    LocalMux I__80 (
            .O(N__768),
            .I(\fsm_shiftRegs_inst1.counterDYNZ0Z_3 ));
    InMux I__79 (
            .O(N__765),
            .I(N__762));
    LocalMux I__78 (
            .O(N__762),
            .I(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3 ));
    InMux I__77 (
            .O(N__759),
            .I(N__755));
    InMux I__76 (
            .O(N__758),
            .I(N__752));
    LocalMux I__75 (
            .O(N__755),
            .I(signal_out_fsm));
    LocalMux I__74 (
            .O(N__752),
            .I(signal_out_fsm));
    InMux I__73 (
            .O(N__747),
            .I(N__744));
    LocalMux I__72 (
            .O(N__744),
            .I(SELSTAT));
    InMux I__71 (
            .O(N__741),
            .I(N__738));
    LocalMux I__70 (
            .O(N__738),
            .I(SELDYN));
    IoInMux I__69 (
            .O(N__735),
            .I(N__732));
    LocalMux I__68 (
            .O(N__732),
            .I(N__729));
    Span12Mux_s0_h I__67 (
            .O(N__729),
            .I(N__726));
    Odrv12 I__66 (
            .O(N__726),
            .I(generated_signal_c));
    IoInMux I__65 (
            .O(N__723),
            .I(N__720));
    LocalMux I__64 (
            .O(N__720),
            .I(RST_N_c_i));
    CascadeMux I__63 (
            .O(N__717),
            .I(\fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_ ));
    defparam IN_MUX_bfv_4_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_11_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB RST_N_ibuf_RNIBJGC_0 (
            .USERSIGNALTOGLOBALBUFFER(N__723),
            .GLOBALBUFFEROUTPUT(RST_N_c_i_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.signal_out_LC_1_10_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.signal_out_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.signal_out_LC_1_10_0 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \fsm_shiftRegs_inst1.signal_out_LC_1_10_0  (
            .in0(N__759),
            .in1(N__906),
            .in2(N__1267),
            .in3(N__1335),
            .lcout(signal_out_fsm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1490),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_RNO_1_2_LC_1_10_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_1_2_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_1_2_LC_1_10_2 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNO_1_2_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__819),
            .in3(N__1039),
            .lcout(\fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.sel_stat_LC_1_11_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.sel_stat_LC_1_11_0 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.sel_stat_LC_1_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fsm_shiftRegs_inst1.sel_stat_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1364),
            .lcout(SELSTAT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1488),
            .ce(),
            .sr(N__1453));
    defparam \fsm_shiftRegs_inst1.sel_dyn_LC_1_11_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.sel_dyn_LC_1_11_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.sel_dyn_LC_1_11_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \fsm_shiftRegs_inst1.sel_dyn_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__1333),
            .in2(_gnd_net_),
            .in3(N__1431),
            .lcout(SELDYN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1488),
            .ce(),
            .sr(N__1453));
    defparam \generator_inst1.signal_aux_LC_1_11_4 .C_ON=1'b0;
    defparam \generator_inst1.signal_aux_LC_1_11_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.signal_aux_LC_1_11_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \generator_inst1.signal_aux_LC_1_11_4  (
            .in0(N__758),
            .in1(N__747),
            .in2(_gnd_net_),
            .in3(N__741),
            .lcout(generated_signal_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1488),
            .ce(),
            .sr(N__1453));
    defparam \fsm_shiftRegs_inst1.current_state_3_LC_1_11_5 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_3_LC_1_11_5 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.current_state_3_LC_1_11_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_3_LC_1_11_5  (
            .in0(N__983),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__765),
            .lcout(\fsm_shiftRegs_inst1.current_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1488),
            .ce(),
            .sr(N__1453));
    defparam RST_N_ibuf_RNIBJGC_LC_1_15_1.C_ON=1'b0;
    defparam RST_N_ibuf_RNIBJGC_LC_1_15_1.SEQ_MODE=4'b0000;
    defparam RST_N_ibuf_RNIBJGC_LC_1_15_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 RST_N_ibuf_RNIBJGC_LC_1_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1268),
            .lcout(RST_N_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_2_LC_2_9_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_2_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_2_LC_2_9_0 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \fsm_shiftRegs_inst1.counter_RNO_0_2_LC_2_9_0  (
            .in0(N__856),
            .in1(N__836),
            .in2(N__1011),
            .in3(N__814),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counter_2_LC_2_9_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_2_LC_2_9_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter_2_LC_2_9_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fsm_shiftRegs_inst1.counter_2_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__717),
            .in3(N__1040),
            .lcout(\fsm_shiftRegs_inst1.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1495),
            .ce(),
            .sr(N__1456));
    defparam \fsm_shiftRegs_inst1.counter_0_LC_2_9_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_0_LC_2_9_2 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter_0_LC_2_9_2 .LUT_INIT=16'b1010000001010000;
    LogicCell40 \fsm_shiftRegs_inst1.counter_0_LC_2_9_2  (
            .in0(N__857),
            .in1(_gnd_net_),
            .in2(N__1047),
            .in3(N__1008),
            .lcout(\fsm_shiftRegs_inst1.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1495),
            .ce(),
            .sr(N__1456));
    defparam \fsm_shiftRegs_inst1.counter_RNIC589_1_LC_2_9_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_RNIC589_1_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.counter_RNIC589_1_LC_2_9_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \fsm_shiftRegs_inst1.counter_RNIC589_1_LC_2_9_3  (
            .in0(N__834),
            .in1(N__854),
            .in2(_gnd_net_),
            .in3(N__1001),
            .lcout(\fsm_shiftRegs_inst1.N_125_1 ),
            .ltout(\fsm_shiftRegs_inst1.N_125_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_1_LC_2_9_4 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_1_LC_2_9_4 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.current_state_1_LC_2_9_4 .LUT_INIT=16'b1110111011001110;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_1_LC_2_9_4  (
            .in0(N__1045),
            .in1(N__1224),
            .in2(N__864),
            .in3(N__815),
            .lcout(\fsm_shiftRegs_inst1.current_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1495),
            .ce(),
            .sr(N__1456));
    defparam \fsm_shiftRegs_inst1.counter_1_LC_2_9_5 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_1_LC_2_9_5 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter_1_LC_2_9_5 .LUT_INIT=16'b1001110000000000;
    LogicCell40 \fsm_shiftRegs_inst1.counter_1_LC_2_9_5  (
            .in0(N__1009),
            .in1(N__837),
            .in2(N__861),
            .in3(N__1044),
            .lcout(\fsm_shiftRegs_inst1.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1495),
            .ce(),
            .sr(N__1456));
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_3_LC_2_9_6 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_3_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.counter_RNO_0_3_LC_2_9_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \fsm_shiftRegs_inst1.counter_RNO_0_3_LC_2_9_6  (
            .in0(N__855),
            .in1(N__835),
            .in2(N__1010),
            .in3(N__813),
            .lcout(\fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counterDYN_RNO_0_3_LC_2_10_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counterDYN_RNO_0_3_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.counterDYN_RNO_0_3_LC_2_10_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \fsm_shiftRegs_inst1.counterDYN_RNO_0_3_LC_2_10_0  (
            .in0(N__950),
            .in1(N__922),
            .in2(N__780),
            .in3(N__976),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counterDYN_3_LC_2_10_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counterDYN_3_LC_2_10_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counterDYN_3_LC_2_10_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fsm_shiftRegs_inst1.counterDYN_3_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__798),
            .in3(N__1331),
            .lcout(\fsm_shiftRegs_inst1.counterDYNZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1493),
            .ce(),
            .sr(N__1454));
    defparam \fsm_shiftRegs_inst1.counterDYN_0_LC_2_10_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counterDYN_0_LC_2_10_2 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counterDYN_0_LC_2_10_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \fsm_shiftRegs_inst1.counterDYN_0_LC_2_10_2  (
            .in0(N__1329),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__980),
            .lcout(\fsm_shiftRegs_inst1.counterDYNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1493),
            .ce(),
            .sr(N__1454));
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_2_LC_2_10_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_2_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_2_LC_2_10_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNO_0_2_LC_2_10_3  (
            .in0(N__923),
            .in1(N__951),
            .in2(N__984),
            .in3(N__779),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_2_LC_2_10_4 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_2_LC_2_10_4 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.current_state_2_LC_2_10_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_2_LC_2_10_4  (
            .in0(N__1330),
            .in1(N__795),
            .in2(N__789),
            .in3(N__786),
            .lcout(\fsm_shiftRegs_inst1.current_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1493),
            .ce(),
            .sr(N__1454));
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_3_LC_2_10_5 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_3_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_3_LC_2_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNO_0_3_LC_2_10_5  (
            .in0(N__921),
            .in1(N__1328),
            .in2(N__954),
            .in3(N__775),
            .lcout(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counterDYN_2_LC_2_10_6 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counterDYN_2_LC_2_10_6 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counterDYN_2_LC_2_10_6 .LUT_INIT=16'b0100100011000000;
    LogicCell40 \fsm_shiftRegs_inst1.counterDYN_2_LC_2_10_6  (
            .in0(N__952),
            .in1(N__1334),
            .in2(N__927),
            .in3(N__981),
            .lcout(\fsm_shiftRegs_inst1.counterDYNZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1493),
            .ce(),
            .sr(N__1454));
    defparam \fsm_shiftRegs_inst1.bit_sequence_15_LC_2_11_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_15_LC_2_11_1 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_15_LC_2_11_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_15_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(N__1212),
            .in2(_gnd_net_),
            .in3(N__900),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1491),
            .ce(N__1286),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_14_LC_2_11_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_14_LC_2_11_2 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_14_LC_2_11_2 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_14_LC_2_11_2  (
            .in0(N__1215),
            .in1(N__894),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1491),
            .ce(N__1286),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_13_LC_2_11_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_13_LC_2_11_3 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_13_LC_2_11_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_13_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__1211),
            .in2(_gnd_net_),
            .in3(N__888),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1491),
            .ce(N__1286),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_12_LC_2_11_4 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_12_LC_2_11_4 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_12_LC_2_11_4 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_12_LC_2_11_4  (
            .in0(N__1214),
            .in1(N__882),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1491),
            .ce(N__1286),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_11_LC_2_11_5 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_11_LC_2_11_5 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_11_LC_2_11_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_11_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__1210),
            .in2(_gnd_net_),
            .in3(N__876),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1491),
            .ce(N__1286),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_10_LC_2_11_6 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_10_LC_2_11_6 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_10_LC_2_11_6 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_10_LC_2_11_6  (
            .in0(N__1213),
            .in1(N__1065),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1491),
            .ce(N__1286),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_6_LC_2_12_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_6_LC_2_12_0 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_6_LC_2_12_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_6_LC_2_12_0  (
            .in0(N__1217),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__870),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1489),
            .ce(N__1287),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_5_LC_2_12_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_5_LC_2_12_1 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_5_LC_2_12_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_5_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__1083),
            .in2(_gnd_net_),
            .in3(N__1220),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1489),
            .ce(N__1287),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_7_LC_2_12_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_7_LC_2_12_2 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_7_LC_2_12_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_7_LC_2_12_2  (
            .in0(N__1218),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1095),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1489),
            .ce(N__1287),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_3_LC_2_12_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_3_LC_2_12_3 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_3_LC_2_12_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_3_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__1154),
            .in2(_gnd_net_),
            .in3(N__1219),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1489),
            .ce(N__1287),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_4_LC_2_12_4 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_4_LC_2_12_4 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_4_LC_2_12_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_4_LC_2_12_4  (
            .in0(N__1216),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1089),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1489),
            .ce(N__1287),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_8_LC_2_12_5 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_8_LC_2_12_5 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_8_LC_2_12_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_8_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(N__1077),
            .in2(_gnd_net_),
            .in3(N__1221),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1489),
            .ce(N__1287),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_9_LC_2_12_7 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_9_LC_2_12_7 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_9_LC_2_12_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_9_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(N__1071),
            .in2(_gnd_net_),
            .in3(N__1222),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1489),
            .ce(N__1287),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.en_fin_LC_2_13_4 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.en_fin_LC_2_13_4 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.en_fin_LC_2_13_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \fsm_shiftRegs_inst1.en_fin_LC_2_13_4  (
            .in0(N__1430),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(ENFIN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1487),
            .ce(),
            .sr(N__1452));
    defparam \fsm_shiftRegs_inst1.counter_3_LC_3_10_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter_3_LC_3_10_0 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter_3_LC_3_10_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fsm_shiftRegs_inst1.counter_3_LC_3_10_0  (
            .in0(_gnd_net_),
            .in1(N__1046),
            .in2(_gnd_net_),
            .in3(N__1017),
            .lcout(\fsm_shiftRegs_inst1.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1496),
            .ce(),
            .sr(N__1457));
    defparam \fsm_shiftRegs_inst1.counterDYN_1_LC_3_10_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counterDYN_1_LC_3_10_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counterDYN_1_LC_3_10_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \fsm_shiftRegs_inst1.counterDYN_1_LC_3_10_1  (
            .in0(N__1332),
            .in1(N__982),
            .in2(_gnd_net_),
            .in3(N__953),
            .lcout(\fsm_shiftRegs_inst1.counterDYNZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1496),
            .ce(),
            .sr(N__1457));
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_4_LC_3_11_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_4_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_4_LC_3_11_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNO_0_4_LC_3_11_0  (
            .in0(N__1116),
            .in1(N__1133),
            .in2(N__1605),
            .in3(N__1568),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_4_LC_3_11_1 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_4_LC_3_11_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.current_state_4_LC_3_11_1 .LUT_INIT=16'b1100111011101110;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_4_LC_3_11_1  (
            .in0(N__1428),
            .in1(N__1365),
            .in2(N__1350),
            .in3(N__1344),
            .lcout(\fsm_shiftRegs_inst1.current_stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1494),
            .ce(),
            .sr(N__1455));
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_0_LC_3_11_2 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_0_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNO_0_0_LC_3_11_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNO_0_0_LC_3_11_2  (
            .in0(N__1601),
            .in1(N__1112),
            .in2(_gnd_net_),
            .in3(N__1567),
            .lcout(),
            .ltout(\fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_0_LC_3_11_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_0_LC_3_11_3 .SEQ_MODE=4'b1011;
    defparam \fsm_shiftRegs_inst1.current_state_0_LC_3_11_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_0_LC_3_11_3  (
            .in0(N__1134),
            .in1(N__1429),
            .in2(N__1347),
            .in3(N__1343),
            .lcout(\fsm_shiftRegs_inst1.current_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1494),
            .ce(),
            .sr(N__1455));
    defparam \fsm_shiftRegs_inst1.counter2_RNITAO81_7_LC_3_11_5 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter2_RNITAO81_7_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.counter2_RNITAO81_7_LC_3_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_RNITAO81_7_LC_3_11_5  (
            .in0(N__1508),
            .in1(N__1583),
            .in2(N__1548),
            .in3(N__1526),
            .lcout(\fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_RNO_0_2_LC_3_11_6 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_RNO_0_2_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_RNO_0_2_LC_3_11_6 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_RNO_0_2_LC_3_11_6  (
            .in0(N__1326),
            .in1(N__1205),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fsm_shiftRegs_inst1.N_122_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.current_state_RNI333L_2_LC_3_11_7 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNI333L_2_LC_3_11_7 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNI333L_2_LC_3_11_7 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNI333L_2_LC_3_11_7  (
            .in0(N__1206),
            .in1(N__1327),
            .in2(_gnd_net_),
            .in3(N__1263),
            .lcout(\fsm_shiftRegs_inst1.un1_current_state4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.bit_sequence_2_LC_3_12_0 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.bit_sequence_2_LC_3_12_0 .SEQ_MODE=4'b1000;
    defparam \fsm_shiftRegs_inst1.bit_sequence_2_LC_3_12_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fsm_shiftRegs_inst1.bit_sequence_2_LC_3_12_0  (
            .in0(N__1269),
            .in1(N__1155),
            .in2(_gnd_net_),
            .in3(N__1223),
            .lcout(\fsm_shiftRegs_inst1.bit_sequenceZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1492),
            .ce(N__1143),
            .sr(_gnd_net_));
    defparam \fsm_shiftRegs_inst1.counter2_0_LC_4_11_0 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_0_LC_4_11_0 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_0_LC_4_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_0_LC_4_11_0  (
            .in0(N__1392),
            .in1(N__1132),
            .in2(_gnd_net_),
            .in3(N__1119),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_0 ),
            .ltout(),
            .carryin(bfn_4_11_0_),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_0 ),
            .clk(N__1497),
            .ce(),
            .sr(N__1458));
    defparam \fsm_shiftRegs_inst1.counter2_1_LC_4_11_1 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_1_LC_4_11_1 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_1_LC_4_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_1_LC_4_11_1  (
            .in0(N__1388),
            .in1(N__1111),
            .in2(_gnd_net_),
            .in3(N__1608),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_1 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_0 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_1 ),
            .clk(N__1497),
            .ce(),
            .sr(N__1458));
    defparam \fsm_shiftRegs_inst1.counter2_2_LC_4_11_2 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_2_LC_4_11_2 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_2_LC_4_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_2_LC_4_11_2  (
            .in0(N__1393),
            .in1(N__1600),
            .in2(_gnd_net_),
            .in3(N__1587),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_2 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_1 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_2 ),
            .clk(N__1497),
            .ce(),
            .sr(N__1458));
    defparam \fsm_shiftRegs_inst1.counter2_3_LC_4_11_3 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_3_LC_4_11_3 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_3_LC_4_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_3_LC_4_11_3  (
            .in0(N__1389),
            .in1(N__1584),
            .in2(_gnd_net_),
            .in3(N__1572),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_3 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_2 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_3 ),
            .clk(N__1497),
            .ce(),
            .sr(N__1458));
    defparam \fsm_shiftRegs_inst1.counter2_4_LC_4_11_4 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_4_LC_4_11_4 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_4_LC_4_11_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_4_LC_4_11_4  (
            .in0(N__1394),
            .in1(_gnd_net_),
            .in2(N__1569),
            .in3(N__1551),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_4 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_3 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_4 ),
            .clk(N__1497),
            .ce(),
            .sr(N__1458));
    defparam \fsm_shiftRegs_inst1.counter2_5_LC_4_11_5 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_5_LC_4_11_5 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_5_LC_4_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_5_LC_4_11_5  (
            .in0(N__1390),
            .in1(N__1547),
            .in2(_gnd_net_),
            .in3(N__1533),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_5 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_4 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_5 ),
            .clk(N__1497),
            .ce(),
            .sr(N__1458));
    defparam \fsm_shiftRegs_inst1.counter2_6_LC_4_11_6 .C_ON=1'b1;
    defparam \fsm_shiftRegs_inst1.counter2_6_LC_4_11_6 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_6_LC_4_11_6 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_6_LC_4_11_6  (
            .in0(N__1395),
            .in1(_gnd_net_),
            .in2(N__1530),
            .in3(N__1515),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_6 ),
            .ltout(),
            .carryin(\fsm_shiftRegs_inst1.counter2_cry_5 ),
            .carryout(\fsm_shiftRegs_inst1.counter2_cry_6 ),
            .clk(N__1497),
            .ce(),
            .sr(N__1458));
    defparam \fsm_shiftRegs_inst1.counter2_7_LC_4_11_7 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.counter2_7_LC_4_11_7 .SEQ_MODE=4'b1010;
    defparam \fsm_shiftRegs_inst1.counter2_7_LC_4_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fsm_shiftRegs_inst1.counter2_7_LC_4_11_7  (
            .in0(N__1391),
            .in1(N__1509),
            .in2(_gnd_net_),
            .in3(N__1512),
            .lcout(\fsm_shiftRegs_inst1.counter2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1497),
            .ce(),
            .sr(N__1458));
    defparam \fsm_shiftRegs_inst1.current_state_RNIVA94_4_LC_4_12_3 .C_ON=1'b0;
    defparam \fsm_shiftRegs_inst1.current_state_RNIVA94_4_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \fsm_shiftRegs_inst1.current_state_RNIVA94_4_LC_4_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \fsm_shiftRegs_inst1.current_state_RNIVA94_4_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1421),
            .lcout(\fsm_shiftRegs_inst1.current_state_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
