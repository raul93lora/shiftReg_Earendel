// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 19 2025 11:24:18

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    SDO_signal_out,
    RST_N,
    CLK_uC,
    CLK);

    output SDO_signal_out;
    input RST_N;
    input CLK_uC;
    input CLK;

    wire N__6294;
    wire N__6293;
    wire N__6292;
    wire N__6283;
    wire N__6282;
    wire N__6281;
    wire N__6274;
    wire N__6273;
    wire N__6272;
    wire N__6265;
    wire N__6264;
    wire N__6263;
    wire N__6246;
    wire N__6243;
    wire N__6240;
    wire N__6237;
    wire N__6234;
    wire N__6231;
    wire N__6228;
    wire N__6225;
    wire N__6222;
    wire N__6219;
    wire N__6216;
    wire N__6213;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6201;
    wire N__6198;
    wire N__6195;
    wire N__6192;
    wire N__6189;
    wire N__6186;
    wire N__6185;
    wire N__6184;
    wire N__6183;
    wire N__6182;
    wire N__6181;
    wire N__6180;
    wire N__6179;
    wire N__6178;
    wire N__6177;
    wire N__6176;
    wire N__6175;
    wire N__6174;
    wire N__6173;
    wire N__6172;
    wire N__6171;
    wire N__6170;
    wire N__6169;
    wire N__6168;
    wire N__6167;
    wire N__6166;
    wire N__6165;
    wire N__6164;
    wire N__6163;
    wire N__6162;
    wire N__6161;
    wire N__6160;
    wire N__6159;
    wire N__6158;
    wire N__6157;
    wire N__6156;
    wire N__6155;
    wire N__6154;
    wire N__6153;
    wire N__6152;
    wire N__6151;
    wire N__6150;
    wire N__6149;
    wire N__6148;
    wire N__6147;
    wire N__6146;
    wire N__6145;
    wire N__6144;
    wire N__6143;
    wire N__6142;
    wire N__6141;
    wire N__6140;
    wire N__6139;
    wire N__6138;
    wire N__6137;
    wire N__6136;
    wire N__6135;
    wire N__6134;
    wire N__6133;
    wire N__6132;
    wire N__6131;
    wire N__6130;
    wire N__6129;
    wire N__6128;
    wire N__6127;
    wire N__6126;
    wire N__6125;
    wire N__6124;
    wire N__6123;
    wire N__6122;
    wire N__6121;
    wire N__6120;
    wire N__6119;
    wire N__5982;
    wire N__5979;
    wire N__5976;
    wire N__5975;
    wire N__5974;
    wire N__5973;
    wire N__5972;
    wire N__5971;
    wire N__5970;
    wire N__5969;
    wire N__5968;
    wire N__5967;
    wire N__5966;
    wire N__5965;
    wire N__5964;
    wire N__5963;
    wire N__5962;
    wire N__5961;
    wire N__5960;
    wire N__5959;
    wire N__5958;
    wire N__5957;
    wire N__5956;
    wire N__5955;
    wire N__5954;
    wire N__5953;
    wire N__5952;
    wire N__5951;
    wire N__5950;
    wire N__5949;
    wire N__5948;
    wire N__5947;
    wire N__5946;
    wire N__5945;
    wire N__5944;
    wire N__5943;
    wire N__5874;
    wire N__5871;
    wire N__5868;
    wire N__5867;
    wire N__5866;
    wire N__5865;
    wire N__5864;
    wire N__5863;
    wire N__5862;
    wire N__5861;
    wire N__5860;
    wire N__5859;
    wire N__5858;
    wire N__5857;
    wire N__5856;
    wire N__5855;
    wire N__5854;
    wire N__5853;
    wire N__5852;
    wire N__5851;
    wire N__5850;
    wire N__5849;
    wire N__5848;
    wire N__5847;
    wire N__5846;
    wire N__5845;
    wire N__5844;
    wire N__5843;
    wire N__5842;
    wire N__5841;
    wire N__5840;
    wire N__5839;
    wire N__5838;
    wire N__5837;
    wire N__5836;
    wire N__5835;
    wire N__5834;
    wire N__5833;
    wire N__5832;
    wire N__5831;
    wire N__5830;
    wire N__5829;
    wire N__5828;
    wire N__5827;
    wire N__5826;
    wire N__5825;
    wire N__5824;
    wire N__5823;
    wire N__5822;
    wire N__5821;
    wire N__5820;
    wire N__5819;
    wire N__5818;
    wire N__5817;
    wire N__5816;
    wire N__5815;
    wire N__5814;
    wire N__5813;
    wire N__5812;
    wire N__5811;
    wire N__5810;
    wire N__5809;
    wire N__5808;
    wire N__5807;
    wire N__5806;
    wire N__5805;
    wire N__5804;
    wire N__5803;
    wire N__5802;
    wire N__5801;
    wire N__5664;
    wire N__5661;
    wire N__5658;
    wire N__5655;
    wire N__5652;
    wire N__5649;
    wire N__5646;
    wire N__5643;
    wire N__5640;
    wire N__5637;
    wire N__5634;
    wire N__5631;
    wire N__5628;
    wire N__5625;
    wire N__5622;
    wire N__5619;
    wire N__5616;
    wire N__5613;
    wire N__5610;
    wire N__5607;
    wire N__5604;
    wire N__5601;
    wire N__5598;
    wire N__5595;
    wire N__5592;
    wire N__5589;
    wire N__5586;
    wire N__5583;
    wire N__5580;
    wire N__5577;
    wire N__5574;
    wire N__5571;
    wire N__5568;
    wire N__5565;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5538;
    wire N__5535;
    wire N__5532;
    wire N__5529;
    wire N__5526;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5514;
    wire N__5511;
    wire N__5508;
    wire N__5505;
    wire N__5502;
    wire N__5499;
    wire N__5496;
    wire N__5493;
    wire N__5490;
    wire N__5487;
    wire N__5484;
    wire N__5481;
    wire N__5478;
    wire N__5475;
    wire N__5472;
    wire N__5469;
    wire N__5466;
    wire N__5463;
    wire N__5460;
    wire N__5457;
    wire N__5454;
    wire N__5451;
    wire N__5448;
    wire N__5445;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5430;
    wire N__5427;
    wire N__5424;
    wire N__5421;
    wire N__5418;
    wire N__5415;
    wire N__5412;
    wire N__5409;
    wire N__5406;
    wire N__5403;
    wire N__5400;
    wire N__5397;
    wire N__5394;
    wire N__5391;
    wire N__5388;
    wire N__5385;
    wire N__5382;
    wire N__5379;
    wire N__5376;
    wire N__5373;
    wire N__5370;
    wire N__5367;
    wire N__5364;
    wire N__5361;
    wire N__5358;
    wire N__5355;
    wire N__5352;
    wire N__5349;
    wire N__5346;
    wire N__5343;
    wire N__5340;
    wire N__5337;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5325;
    wire N__5322;
    wire N__5319;
    wire N__5316;
    wire N__5313;
    wire N__5310;
    wire N__5307;
    wire N__5304;
    wire N__5301;
    wire N__5298;
    wire N__5295;
    wire N__5292;
    wire N__5289;
    wire N__5286;
    wire N__5283;
    wire N__5280;
    wire N__5277;
    wire N__5274;
    wire N__5271;
    wire N__5268;
    wire N__5265;
    wire N__5262;
    wire N__5259;
    wire N__5256;
    wire N__5253;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5208;
    wire N__5205;
    wire N__5202;
    wire N__5199;
    wire N__5196;
    wire N__5193;
    wire N__5190;
    wire N__5187;
    wire N__5184;
    wire N__5181;
    wire N__5178;
    wire N__5175;
    wire N__5172;
    wire N__5169;
    wire N__5166;
    wire N__5163;
    wire N__5160;
    wire N__5157;
    wire N__5154;
    wire N__5153;
    wire N__5152;
    wire N__5149;
    wire N__5146;
    wire N__5145;
    wire N__5142;
    wire N__5137;
    wire N__5134;
    wire N__5131;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5115;
    wire N__5114;
    wire N__5113;
    wire N__5112;
    wire N__5109;
    wire N__5106;
    wire N__5099;
    wire N__5094;
    wire N__5093;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5076;
    wire N__5075;
    wire N__5074;
    wire N__5073;
    wire N__5070;
    wire N__5063;
    wire N__5060;
    wire N__5055;
    wire N__5054;
    wire N__5053;
    wire N__5052;
    wire N__5051;
    wire N__5050;
    wire N__5049;
    wire N__5048;
    wire N__5047;
    wire N__5046;
    wire N__5045;
    wire N__5040;
    wire N__5039;
    wire N__5038;
    wire N__5037;
    wire N__5036;
    wire N__5025;
    wire N__5024;
    wire N__5023;
    wire N__5022;
    wire N__5019;
    wire N__5012;
    wire N__5011;
    wire N__5010;
    wire N__5009;
    wire N__5008;
    wire N__5007;
    wire N__5006;
    wire N__5005;
    wire N__5004;
    wire N__5003;
    wire N__5002;
    wire N__5001;
    wire N__5000;
    wire N__4999;
    wire N__4998;
    wire N__4997;
    wire N__4996;
    wire N__4995;
    wire N__4994;
    wire N__4993;
    wire N__4992;
    wire N__4991;
    wire N__4990;
    wire N__4989;
    wire N__4988;
    wire N__4987;
    wire N__4986;
    wire N__4985;
    wire N__4984;
    wire N__4983;
    wire N__4980;
    wire N__4973;
    wire N__4972;
    wire N__4971;
    wire N__4970;
    wire N__4969;
    wire N__4968;
    wire N__4967;
    wire N__4966;
    wire N__4965;
    wire N__4964;
    wire N__4963;
    wire N__4962;
    wire N__4961;
    wire N__4960;
    wire N__4957;
    wire N__4956;
    wire N__4955;
    wire N__4954;
    wire N__4953;
    wire N__4952;
    wire N__4951;
    wire N__4950;
    wire N__4949;
    wire N__4948;
    wire N__4947;
    wire N__4946;
    wire N__4945;
    wire N__4944;
    wire N__4943;
    wire N__4942;
    wire N__4939;
    wire N__4932;
    wire N__4927;
    wire N__4922;
    wire N__4911;
    wire N__4900;
    wire N__4885;
    wire N__4868;
    wire N__4867;
    wire N__4866;
    wire N__4865;
    wire N__4864;
    wire N__4863;
    wire N__4862;
    wire N__4861;
    wire N__4860;
    wire N__4859;
    wire N__4858;
    wire N__4857;
    wire N__4856;
    wire N__4855;
    wire N__4854;
    wire N__4853;
    wire N__4852;
    wire N__4847;
    wire N__4842;
    wire N__4839;
    wire N__4828;
    wire N__4823;
    wire N__4814;
    wire N__4811;
    wire N__4810;
    wire N__4809;
    wire N__4808;
    wire N__4807;
    wire N__4806;
    wire N__4803;
    wire N__4788;
    wire N__4771;
    wire N__4756;
    wire N__4753;
    wire N__4738;
    wire N__4721;
    wire N__4718;
    wire N__4707;
    wire N__4704;
    wire N__4701;
    wire N__4698;
    wire N__4695;
    wire N__4694;
    wire N__4691;
    wire N__4690;
    wire N__4689;
    wire N__4688;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4674;
    wire N__4665;
    wire N__4656;
    wire N__4651;
    wire N__4648;
    wire N__4643;
    wire N__4636;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4596;
    wire N__4595;
    wire N__4594;
    wire N__4593;
    wire N__4592;
    wire N__4591;
    wire N__4590;
    wire N__4589;
    wire N__4588;
    wire N__4585;
    wire N__4584;
    wire N__4583;
    wire N__4570;
    wire N__4569;
    wire N__4568;
    wire N__4567;
    wire N__4566;
    wire N__4565;
    wire N__4560;
    wire N__4557;
    wire N__4556;
    wire N__4555;
    wire N__4554;
    wire N__4553;
    wire N__4552;
    wire N__4551;
    wire N__4550;
    wire N__4549;
    wire N__4548;
    wire N__4547;
    wire N__4546;
    wire N__4545;
    wire N__4544;
    wire N__4543;
    wire N__4542;
    wire N__4541;
    wire N__4536;
    wire N__4533;
    wire N__4522;
    wire N__4517;
    wire N__4510;
    wire N__4509;
    wire N__4508;
    wire N__4507;
    wire N__4504;
    wire N__4487;
    wire N__4482;
    wire N__4477;
    wire N__4466;
    wire N__4459;
    wire N__4446;
    wire N__4443;
    wire N__4442;
    wire N__4441;
    wire N__4440;
    wire N__4439;
    wire N__4436;
    wire N__4429;
    wire N__4426;
    wire N__4419;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4404;
    wire N__4401;
    wire N__4398;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4368;
    wire N__4365;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4328;
    wire N__4327;
    wire N__4326;
    wire N__4317;
    wire N__4314;
    wire N__4313;
    wire N__4312;
    wire N__4309;
    wire N__4306;
    wire N__4303;
    wire N__4296;
    wire N__4293;
    wire N__4292;
    wire N__4289;
    wire N__4288;
    wire N__4287;
    wire N__4286;
    wire N__4275;
    wire N__4272;
    wire N__4271;
    wire N__4270;
    wire N__4269;
    wire N__4268;
    wire N__4267;
    wire N__4264;
    wire N__4255;
    wire N__4252;
    wire N__4247;
    wire N__4242;
    wire N__4239;
    wire N__4236;
    wire N__4233;
    wire N__4230;
    wire N__4227;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4217;
    wire N__4216;
    wire N__4215;
    wire N__4214;
    wire N__4213;
    wire N__4212;
    wire N__4211;
    wire N__4210;
    wire N__4209;
    wire N__4208;
    wire N__4207;
    wire N__4206;
    wire N__4205;
    wire N__4204;
    wire N__4203;
    wire N__4202;
    wire N__4201;
    wire N__4200;
    wire N__4199;
    wire N__4198;
    wire N__4155;
    wire N__4152;
    wire N__4149;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4128;
    wire N__4125;
    wire N__4122;
    wire N__4121;
    wire N__4120;
    wire N__4119;
    wire N__4118;
    wire N__4117;
    wire N__4116;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4086;
    wire N__4085;
    wire N__4084;
    wire N__4081;
    wire N__4078;
    wire N__4077;
    wire N__4076;
    wire N__4075;
    wire N__4074;
    wire N__4071;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4044;
    wire N__4043;
    wire N__4042;
    wire N__4039;
    wire N__4036;
    wire N__4033;
    wire N__4026;
    wire N__4023;
    wire N__4020;
    wire N__4017;
    wire N__4014;
    wire N__4013;
    wire N__4012;
    wire N__4011;
    wire N__4010;
    wire N__4007;
    wire N__4006;
    wire N__4005;
    wire N__4002;
    wire N__3999;
    wire N__3996;
    wire N__3993;
    wire N__3990;
    wire N__3983;
    wire N__3972;
    wire N__3971;
    wire N__3970;
    wire N__3969;
    wire N__3968;
    wire N__3967;
    wire N__3966;
    wire N__3963;
    wire N__3958;
    wire N__3955;
    wire N__3950;
    wire N__3947;
    wire N__3936;
    wire N__3933;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3921;
    wire N__3918;
    wire N__3915;
    wire N__3912;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3900;
    wire N__3897;
    wire N__3894;
    wire N__3891;
    wire N__3888;
    wire N__3885;
    wire N__3882;
    wire N__3879;
    wire N__3876;
    wire N__3873;
    wire N__3870;
    wire N__3867;
    wire N__3864;
    wire N__3861;
    wire N__3858;
    wire N__3855;
    wire N__3852;
    wire N__3849;
    wire N__3846;
    wire N__3843;
    wire N__3840;
    wire N__3837;
    wire N__3834;
    wire N__3831;
    wire N__3828;
    wire N__3825;
    wire N__3822;
    wire N__3819;
    wire N__3816;
    wire N__3813;
    wire N__3810;
    wire N__3807;
    wire N__3804;
    wire N__3801;
    wire N__3798;
    wire N__3795;
    wire N__3792;
    wire N__3789;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3771;
    wire N__3768;
    wire N__3765;
    wire N__3762;
    wire N__3759;
    wire N__3756;
    wire N__3753;
    wire N__3750;
    wire N__3747;
    wire N__3744;
    wire N__3741;
    wire N__3738;
    wire N__3735;
    wire N__3732;
    wire N__3729;
    wire N__3726;
    wire N__3723;
    wire N__3720;
    wire N__3717;
    wire N__3714;
    wire N__3711;
    wire N__3708;
    wire N__3705;
    wire N__3702;
    wire N__3699;
    wire N__3696;
    wire N__3693;
    wire N__3690;
    wire N__3687;
    wire N__3684;
    wire N__3681;
    wire N__3678;
    wire N__3675;
    wire N__3672;
    wire N__3669;
    wire N__3666;
    wire N__3663;
    wire N__3660;
    wire N__3657;
    wire N__3654;
    wire N__3651;
    wire N__3648;
    wire N__3645;
    wire N__3642;
    wire N__3639;
    wire N__3638;
    wire N__3637;
    wire N__3636;
    wire N__3631;
    wire N__3626;
    wire N__3621;
    wire N__3618;
    wire N__3615;
    wire N__3612;
    wire N__3609;
    wire N__3606;
    wire N__3603;
    wire N__3600;
    wire N__3597;
    wire N__3594;
    wire N__3591;
    wire N__3588;
    wire N__3585;
    wire N__3582;
    wire N__3579;
    wire N__3576;
    wire N__3573;
    wire N__3570;
    wire N__3567;
    wire N__3564;
    wire N__3561;
    wire N__3558;
    wire N__3555;
    wire N__3552;
    wire N__3549;
    wire N__3546;
    wire N__3543;
    wire N__3540;
    wire N__3537;
    wire N__3534;
    wire N__3531;
    wire N__3528;
    wire N__3525;
    wire N__3522;
    wire N__3519;
    wire N__3516;
    wire N__3513;
    wire N__3510;
    wire N__3507;
    wire N__3504;
    wire N__3501;
    wire N__3498;
    wire N__3495;
    wire N__3492;
    wire N__3489;
    wire N__3486;
    wire N__3483;
    wire N__3480;
    wire N__3477;
    wire N__3474;
    wire N__3471;
    wire N__3468;
    wire N__3465;
    wire N__3462;
    wire N__3459;
    wire N__3456;
    wire N__3453;
    wire N__3450;
    wire N__3447;
    wire N__3444;
    wire N__3441;
    wire N__3438;
    wire N__3435;
    wire N__3432;
    wire N__3429;
    wire N__3426;
    wire N__3423;
    wire N__3420;
    wire N__3417;
    wire N__3414;
    wire N__3411;
    wire N__3408;
    wire N__3405;
    wire N__3402;
    wire N__3399;
    wire N__3396;
    wire N__3393;
    wire N__3390;
    wire N__3387;
    wire N__3384;
    wire N__3381;
    wire N__3378;
    wire N__3375;
    wire N__3372;
    wire N__3369;
    wire N__3366;
    wire N__3363;
    wire N__3360;
    wire N__3357;
    wire N__3354;
    wire N__3351;
    wire N__3348;
    wire N__3345;
    wire N__3342;
    wire N__3339;
    wire N__3336;
    wire N__3333;
    wire N__3330;
    wire N__3327;
    wire N__3326;
    wire N__3325;
    wire N__3322;
    wire N__3319;
    wire N__3316;
    wire N__3313;
    wire N__3308;
    wire N__3303;
    wire N__3300;
    wire N__3297;
    wire N__3294;
    wire N__3291;
    wire N__3288;
    wire N__3285;
    wire N__3282;
    wire N__3279;
    wire N__3276;
    wire N__3273;
    wire N__3270;
    wire N__3267;
    wire N__3264;
    wire N__3261;
    wire N__3258;
    wire N__3255;
    wire N__3252;
    wire N__3249;
    wire N__3246;
    wire N__3243;
    wire N__3240;
    wire N__3237;
    wire N__3234;
    wire N__3231;
    wire N__3228;
    wire N__3225;
    wire N__3222;
    wire N__3219;
    wire N__3216;
    wire N__3213;
    wire N__3210;
    wire N__3207;
    wire N__3204;
    wire N__3201;
    wire N__3198;
    wire N__3195;
    wire N__3192;
    wire N__3189;
    wire N__3186;
    wire N__3183;
    wire N__3180;
    wire N__3177;
    wire N__3174;
    wire N__3171;
    wire N__3168;
    wire N__3165;
    wire N__3162;
    wire N__3159;
    wire N__3156;
    wire N__3153;
    wire N__3150;
    wire N__3147;
    wire N__3144;
    wire N__3141;
    wire N__3138;
    wire N__3135;
    wire N__3132;
    wire VCCG0;
    wire GNDG0;
    wire RST_N_c;
    wire RST_N_c_i;
    wire \fsm_ctrl_inst1.current_state_i_0 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_58 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_57 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_6 ;
    wire \fsm_ctrl_inst1.bit_sequence_dinZ0Z_0 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_84 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_85 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_86 ;
    wire \fsm_ctrl_inst1.bit_sequence_dinZ0Z_1 ;
    wire \fsm_ctrl_inst1.bit_sequence_dinZ0Z_2 ;
    wire \fsm_ctrl_inst1.bit_sequence_dinZ0Z_5 ;
    wire \fsm_ctrl_inst1.bit_sequence_dinZ0Z_3 ;
    wire \fsm_ctrl_inst1.bit_sequence_dinZ0Z_4 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_56 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_59 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_55 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_7 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_8 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_9 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_10 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_83 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_42 ;
    wire bfn_3_20_0_;
    wire \fsm_ctrl_inst1.counter_idle_cry_0 ;
    wire \fsm_ctrl_inst1.counter_idle_cry_1 ;
    wire \fsm_ctrl_inst1.counter_idle_cry_2 ;
    wire \fsm_ctrl_inst1.counter_idle_cry_3 ;
    wire \fsm_ctrl_inst1.bit_sequence_dinZ0Z_9 ;
    wire \fsm_ctrl_inst1.bit_sequence_dinZ0Z_6 ;
    wire \fsm_ctrl_inst1.bit_sequence_dinZ0Z_7 ;
    wire \fsm_ctrl_inst1.bit_sequence_dinZ0Z_8 ;
    wire \fsm_ctrl_inst1.bit_sequence_dinZ0Z_12 ;
    wire \fsm_ctrl_inst1.bit_sequence_dinZ0Z_10 ;
    wire \fsm_ctrl_inst1.bit_sequence_dinZ0Z_11 ;
    wire \fsm_ctrl_inst1.bit_sequence_dinZ0Z_13 ;
    wire \fsm_ctrl_inst1.bit_sequence_dinZ0Z_14 ;
    wire \fsm_ctrl_inst1.current_state_i_1 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_75 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_76 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_77 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_11 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_54 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_60 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_61 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_78 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_79 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_80 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_4 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_5 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_53 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_37 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_81 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_82 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_3 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_1 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_2 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_38 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_39 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_0 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_40 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_41 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_43 ;
    wire \fsm_ctrl_inst1.g0_0_2_0_cascade_ ;
    wire \fsm_ctrl_inst1.counter_idle_s_3 ;
    wire \fsm_ctrl_inst1.g0_0_2_cascade_ ;
    wire \fsm_ctrl_inst1.counter_idle_s_4 ;
    wire \fsm_ctrl_inst1.g0_0_3_1 ;
    wire \fsm_ctrl_inst1.g0_0_2_1 ;
    wire \fsm_ctrl_inst1.current_state_20_d_i_cascade_ ;
    wire \fsm_ctrl_inst1.counter_idle_s_2 ;
    wire \fsm_ctrl_inst1.N_93_0_cascade_ ;
    wire \fsm_ctrl_inst1.counter_idle_RNO_1Z0Z_0_cascade_ ;
    wire \fsm_ctrl_inst1.counter_idlee_0_cascade_ ;
    wire \fsm_ctrl_inst1.counter_idle_s_1 ;
    wire \fsm_ctrl_inst1.g0_0_3_2 ;
    wire \fsm_ctrl_inst1.g0_0_2_2 ;
    wire \fsm_ctrl_inst1.current_state_20_d_i ;
    wire \fsm_ctrl_inst1.bit_sequence_dinZ0Z_15 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_87 ;
    wire CONSTANT_ONE_NET;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_67 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_64 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_65 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_66 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_68 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_69 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_70 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_73 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_74 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_71 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_72 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_18 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_17 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_16 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_14 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_15 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_62 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_63 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_21 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_22 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_48 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_26 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_12 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_13 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_49 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_50 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_47 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_25 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_44 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_51 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_52 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_23 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_24 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_45 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_46 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_27 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_28 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_33 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_29 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_34 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_30 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_35 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_36 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_31 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_32 ;
    wire \fsm_ctrl_inst1.counter_idleZ0Z_1 ;
    wire \fsm_ctrl_inst1.counter_idleZ0Z_3 ;
    wire \fsm_ctrl_inst1.counter_idleZ0Z_0 ;
    wire \fsm_ctrl_inst1.current_state_RNO_2Z0Z_0 ;
    wire \fsm_ctrl_inst1.g0_0_3_0 ;
    wire \fsm_ctrl_inst1.counter_idleZ1Z_4 ;
    wire \fsm_ctrl_inst1.counter_idleZ0Z_2 ;
    wire \fsm_ctrl_inst1.g0_0_3 ;
    wire \fsm_ctrl_inst1.counter_din_RNO_0Z0Z_3_cascade_ ;
    wire \fsm_ctrl_inst1.current_state_RNO_3Z0Z_0_cascade_ ;
    wire \fsm_ctrl_inst1.current_state_RNO_1Z0Z_0 ;
    wire \fsm_ctrl_inst1.counter_dinZ0Z_2 ;
    wire \fsm_ctrl_inst1.counter_dinZ0Z_3 ;
    wire \fsm_ctrl_inst1.counter_dinZ0Z_1 ;
    wire \fsm_ctrl_inst1.counter_dinZ0Z_0 ;
    wire \fsm_ctrl_inst1.o2_cascade_ ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_0 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_19 ;
    wire \fsm_ctrl_inst1.bit_sequence_statZ0Z_20 ;
    wire \fsm_ctrl_inst1.current_state_i_g_0 ;
    wire SDO_signal_out_c;
    wire \config_register_latched_dec_inst1.DYNSRZ0Z_14 ;
    wire \config_register_latched_dec_inst1.DYNSRZ0Z_15 ;
    wire \config_register_latched_dec_inst1.DYNSRZ0Z_12 ;
    wire \config_register_latched_dec_inst1.DYNSRZ0Z_13 ;
    wire \config_register_latched_dec_inst1.DYNSRZ0Z_10 ;
    wire \config_register_latched_dec_inst1.DYNSRZ0Z_11 ;
    wire \config_register_latched_dec_inst1.DYNSR_cnv_x0Z0Z_0_cascade_ ;
    wire \config_register_latched_dec_inst1.DYNSR_cnv_x1Z0Z_0 ;
    wire CLK_uC_c;
    wire fsm_ctrl_inst1_SCLK_i;
    wire fsm_ctrl_inst1_current_state_1;
    wire \config_register_latched_dec_inst1.STATSR_cnv_x1Z0Z_0_cascade_ ;
    wire \config_register_latched_dec_inst1.STATSR_cnv_x0Z0Z_0 ;
    wire STATSR_cnv_ns_0;
    wire fsm_ctrl_inst1_current_state_0;
    wire SEL_REG;
    wire MOSI;
    wire \config_register_latched_dec_inst1.DYNSRZ0Z_0 ;
    wire \config_register_latched_dec_inst1.DYNSRZ0Z_1 ;
    wire \config_register_latched_dec_inst1.DYNSRZ0Z_2 ;
    wire \config_register_latched_dec_inst1.DYNSRZ0Z_3 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_1 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_2 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_3 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_87 ;
    wire \config_register_latched_dec_inst1.DYNSRZ0Z_9 ;
    wire \config_register_latched_dec_inst1.DYNSRZ0Z_6 ;
    wire \config_register_latched_dec_inst1.DYNSRZ0Z_7 ;
    wire \config_register_latched_dec_inst1.DYNSRZ0Z_8 ;
    wire \config_register_latched_dec_inst1.DYNSRZ0Z_4 ;
    wire \config_register_latched_dec_inst1.DYNSRZ0Z_5 ;
    wire \config_register_latched_dec_inst1.DYNSR_cnv_nsZ0Z_0 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_4 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_5 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_86 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_6 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_7 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_8 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_84 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_85 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_9 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_10 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_11 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_83 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_12 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_81 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_82 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_13 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_80 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_79 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_77 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_78 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_14 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_75 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_76 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_74 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_15 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_16 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_73 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_17 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_18 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_71 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_72 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_70 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_68 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_69 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_67 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_66 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_19 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_20 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_41 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_40 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_42 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_43 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_44 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_45 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_21 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_65 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_36 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_35 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_37 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_38 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_39 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_46 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_47 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_22 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_48 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_23 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_49 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_52 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_50 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_51 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_64 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_63 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_53 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_61 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_62 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_30 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_34 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_31 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_32 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_33 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_26 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_24 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_25 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_27 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_28 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_29 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_60 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_54 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_59 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_57 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_58 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_55 ;
    wire \config_register_latched_dec_inst1.STATSRZ0Z_56 ;
    wire _gnd_net_;
    wire CLK_0_c_g;
    wire N_218_g;
    wire RST_N_c_i_g;

    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6292),
            .GLOBALBUFFEROUTPUT(CLK_0_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__6294),
            .DIN(N__6293),
            .DOUT(N__6292),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__6294),
            .PADOUT(N__6293),
            .PADIN(N__6292),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_uC_ibuf_iopad (
            .OE(N__6283),
            .DIN(N__6282),
            .DOUT(N__6281),
            .PACKAGEPIN(CLK_uC));
    defparam CLK_uC_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_uC_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_uC_ibuf_preio (
            .PADOEN(N__6283),
            .PADOUT(N__6282),
            .PADIN(N__6281),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK_uC_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RST_N_ibuf_iopad (
            .OE(N__6274),
            .DIN(N__6273),
            .DOUT(N__6272),
            .PACKAGEPIN(RST_N));
    defparam RST_N_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RST_N_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RST_N_ibuf_preio (
            .PADOEN(N__6274),
            .PADOUT(N__6273),
            .PADIN(N__6272),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RST_N_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SDO_signal_out_obuf_iopad (
            .OE(N__6265),
            .DIN(N__6264),
            .DOUT(N__6263),
            .PACKAGEPIN(SDO_signal_out));
    defparam SDO_signal_out_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SDO_signal_out_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SDO_signal_out_obuf_preio (
            .PADOEN(N__6265),
            .PADOUT(N__6264),
            .PADIN(N__6263),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4149),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1304 (
            .O(N__6246),
            .I(N__6243));
    LocalMux I__1303 (
            .O(N__6243),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_27 ));
    InMux I__1302 (
            .O(N__6240),
            .I(N__6237));
    LocalMux I__1301 (
            .O(N__6237),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_28 ));
    InMux I__1300 (
            .O(N__6234),
            .I(N__6231));
    LocalMux I__1299 (
            .O(N__6231),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_29 ));
    InMux I__1298 (
            .O(N__6228),
            .I(N__6225));
    LocalMux I__1297 (
            .O(N__6225),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_60 ));
    InMux I__1296 (
            .O(N__6222),
            .I(N__6219));
    LocalMux I__1295 (
            .O(N__6219),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_54 ));
    InMux I__1294 (
            .O(N__6216),
            .I(N__6213));
    LocalMux I__1293 (
            .O(N__6213),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_59 ));
    InMux I__1292 (
            .O(N__6210),
            .I(N__6207));
    LocalMux I__1291 (
            .O(N__6207),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_57 ));
    InMux I__1290 (
            .O(N__6204),
            .I(N__6201));
    LocalMux I__1289 (
            .O(N__6201),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_58 ));
    InMux I__1288 (
            .O(N__6198),
            .I(N__6195));
    LocalMux I__1287 (
            .O(N__6195),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_55 ));
    InMux I__1286 (
            .O(N__6192),
            .I(N__6189));
    LocalMux I__1285 (
            .O(N__6189),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_56 ));
    ClkMux I__1284 (
            .O(N__6186),
            .I(N__5982));
    ClkMux I__1283 (
            .O(N__6185),
            .I(N__5982));
    ClkMux I__1282 (
            .O(N__6184),
            .I(N__5982));
    ClkMux I__1281 (
            .O(N__6183),
            .I(N__5982));
    ClkMux I__1280 (
            .O(N__6182),
            .I(N__5982));
    ClkMux I__1279 (
            .O(N__6181),
            .I(N__5982));
    ClkMux I__1278 (
            .O(N__6180),
            .I(N__5982));
    ClkMux I__1277 (
            .O(N__6179),
            .I(N__5982));
    ClkMux I__1276 (
            .O(N__6178),
            .I(N__5982));
    ClkMux I__1275 (
            .O(N__6177),
            .I(N__5982));
    ClkMux I__1274 (
            .O(N__6176),
            .I(N__5982));
    ClkMux I__1273 (
            .O(N__6175),
            .I(N__5982));
    ClkMux I__1272 (
            .O(N__6174),
            .I(N__5982));
    ClkMux I__1271 (
            .O(N__6173),
            .I(N__5982));
    ClkMux I__1270 (
            .O(N__6172),
            .I(N__5982));
    ClkMux I__1269 (
            .O(N__6171),
            .I(N__5982));
    ClkMux I__1268 (
            .O(N__6170),
            .I(N__5982));
    ClkMux I__1267 (
            .O(N__6169),
            .I(N__5982));
    ClkMux I__1266 (
            .O(N__6168),
            .I(N__5982));
    ClkMux I__1265 (
            .O(N__6167),
            .I(N__5982));
    ClkMux I__1264 (
            .O(N__6166),
            .I(N__5982));
    ClkMux I__1263 (
            .O(N__6165),
            .I(N__5982));
    ClkMux I__1262 (
            .O(N__6164),
            .I(N__5982));
    ClkMux I__1261 (
            .O(N__6163),
            .I(N__5982));
    ClkMux I__1260 (
            .O(N__6162),
            .I(N__5982));
    ClkMux I__1259 (
            .O(N__6161),
            .I(N__5982));
    ClkMux I__1258 (
            .O(N__6160),
            .I(N__5982));
    ClkMux I__1257 (
            .O(N__6159),
            .I(N__5982));
    ClkMux I__1256 (
            .O(N__6158),
            .I(N__5982));
    ClkMux I__1255 (
            .O(N__6157),
            .I(N__5982));
    ClkMux I__1254 (
            .O(N__6156),
            .I(N__5982));
    ClkMux I__1253 (
            .O(N__6155),
            .I(N__5982));
    ClkMux I__1252 (
            .O(N__6154),
            .I(N__5982));
    ClkMux I__1251 (
            .O(N__6153),
            .I(N__5982));
    ClkMux I__1250 (
            .O(N__6152),
            .I(N__5982));
    ClkMux I__1249 (
            .O(N__6151),
            .I(N__5982));
    ClkMux I__1248 (
            .O(N__6150),
            .I(N__5982));
    ClkMux I__1247 (
            .O(N__6149),
            .I(N__5982));
    ClkMux I__1246 (
            .O(N__6148),
            .I(N__5982));
    ClkMux I__1245 (
            .O(N__6147),
            .I(N__5982));
    ClkMux I__1244 (
            .O(N__6146),
            .I(N__5982));
    ClkMux I__1243 (
            .O(N__6145),
            .I(N__5982));
    ClkMux I__1242 (
            .O(N__6144),
            .I(N__5982));
    ClkMux I__1241 (
            .O(N__6143),
            .I(N__5982));
    ClkMux I__1240 (
            .O(N__6142),
            .I(N__5982));
    ClkMux I__1239 (
            .O(N__6141),
            .I(N__5982));
    ClkMux I__1238 (
            .O(N__6140),
            .I(N__5982));
    ClkMux I__1237 (
            .O(N__6139),
            .I(N__5982));
    ClkMux I__1236 (
            .O(N__6138),
            .I(N__5982));
    ClkMux I__1235 (
            .O(N__6137),
            .I(N__5982));
    ClkMux I__1234 (
            .O(N__6136),
            .I(N__5982));
    ClkMux I__1233 (
            .O(N__6135),
            .I(N__5982));
    ClkMux I__1232 (
            .O(N__6134),
            .I(N__5982));
    ClkMux I__1231 (
            .O(N__6133),
            .I(N__5982));
    ClkMux I__1230 (
            .O(N__6132),
            .I(N__5982));
    ClkMux I__1229 (
            .O(N__6131),
            .I(N__5982));
    ClkMux I__1228 (
            .O(N__6130),
            .I(N__5982));
    ClkMux I__1227 (
            .O(N__6129),
            .I(N__5982));
    ClkMux I__1226 (
            .O(N__6128),
            .I(N__5982));
    ClkMux I__1225 (
            .O(N__6127),
            .I(N__5982));
    ClkMux I__1224 (
            .O(N__6126),
            .I(N__5982));
    ClkMux I__1223 (
            .O(N__6125),
            .I(N__5982));
    ClkMux I__1222 (
            .O(N__6124),
            .I(N__5982));
    ClkMux I__1221 (
            .O(N__6123),
            .I(N__5982));
    ClkMux I__1220 (
            .O(N__6122),
            .I(N__5982));
    ClkMux I__1219 (
            .O(N__6121),
            .I(N__5982));
    ClkMux I__1218 (
            .O(N__6120),
            .I(N__5982));
    ClkMux I__1217 (
            .O(N__6119),
            .I(N__5982));
    GlobalMux I__1216 (
            .O(N__5982),
            .I(N__5979));
    gio2CtrlBuf I__1215 (
            .O(N__5979),
            .I(CLK_0_c_g));
    CEMux I__1214 (
            .O(N__5976),
            .I(N__5874));
    CEMux I__1213 (
            .O(N__5975),
            .I(N__5874));
    CEMux I__1212 (
            .O(N__5974),
            .I(N__5874));
    CEMux I__1211 (
            .O(N__5973),
            .I(N__5874));
    CEMux I__1210 (
            .O(N__5972),
            .I(N__5874));
    CEMux I__1209 (
            .O(N__5971),
            .I(N__5874));
    CEMux I__1208 (
            .O(N__5970),
            .I(N__5874));
    CEMux I__1207 (
            .O(N__5969),
            .I(N__5874));
    CEMux I__1206 (
            .O(N__5968),
            .I(N__5874));
    CEMux I__1205 (
            .O(N__5967),
            .I(N__5874));
    CEMux I__1204 (
            .O(N__5966),
            .I(N__5874));
    CEMux I__1203 (
            .O(N__5965),
            .I(N__5874));
    CEMux I__1202 (
            .O(N__5964),
            .I(N__5874));
    CEMux I__1201 (
            .O(N__5963),
            .I(N__5874));
    CEMux I__1200 (
            .O(N__5962),
            .I(N__5874));
    CEMux I__1199 (
            .O(N__5961),
            .I(N__5874));
    CEMux I__1198 (
            .O(N__5960),
            .I(N__5874));
    CEMux I__1197 (
            .O(N__5959),
            .I(N__5874));
    CEMux I__1196 (
            .O(N__5958),
            .I(N__5874));
    CEMux I__1195 (
            .O(N__5957),
            .I(N__5874));
    CEMux I__1194 (
            .O(N__5956),
            .I(N__5874));
    CEMux I__1193 (
            .O(N__5955),
            .I(N__5874));
    CEMux I__1192 (
            .O(N__5954),
            .I(N__5874));
    CEMux I__1191 (
            .O(N__5953),
            .I(N__5874));
    CEMux I__1190 (
            .O(N__5952),
            .I(N__5874));
    CEMux I__1189 (
            .O(N__5951),
            .I(N__5874));
    CEMux I__1188 (
            .O(N__5950),
            .I(N__5874));
    CEMux I__1187 (
            .O(N__5949),
            .I(N__5874));
    CEMux I__1186 (
            .O(N__5948),
            .I(N__5874));
    CEMux I__1185 (
            .O(N__5947),
            .I(N__5874));
    CEMux I__1184 (
            .O(N__5946),
            .I(N__5874));
    CEMux I__1183 (
            .O(N__5945),
            .I(N__5874));
    CEMux I__1182 (
            .O(N__5944),
            .I(N__5874));
    CEMux I__1181 (
            .O(N__5943),
            .I(N__5874));
    GlobalMux I__1180 (
            .O(N__5874),
            .I(N__5871));
    gio2CtrlBuf I__1179 (
            .O(N__5871),
            .I(N_218_g));
    SRMux I__1178 (
            .O(N__5868),
            .I(N__5664));
    SRMux I__1177 (
            .O(N__5867),
            .I(N__5664));
    SRMux I__1176 (
            .O(N__5866),
            .I(N__5664));
    SRMux I__1175 (
            .O(N__5865),
            .I(N__5664));
    SRMux I__1174 (
            .O(N__5864),
            .I(N__5664));
    SRMux I__1173 (
            .O(N__5863),
            .I(N__5664));
    SRMux I__1172 (
            .O(N__5862),
            .I(N__5664));
    SRMux I__1171 (
            .O(N__5861),
            .I(N__5664));
    SRMux I__1170 (
            .O(N__5860),
            .I(N__5664));
    SRMux I__1169 (
            .O(N__5859),
            .I(N__5664));
    SRMux I__1168 (
            .O(N__5858),
            .I(N__5664));
    SRMux I__1167 (
            .O(N__5857),
            .I(N__5664));
    SRMux I__1166 (
            .O(N__5856),
            .I(N__5664));
    SRMux I__1165 (
            .O(N__5855),
            .I(N__5664));
    SRMux I__1164 (
            .O(N__5854),
            .I(N__5664));
    SRMux I__1163 (
            .O(N__5853),
            .I(N__5664));
    SRMux I__1162 (
            .O(N__5852),
            .I(N__5664));
    SRMux I__1161 (
            .O(N__5851),
            .I(N__5664));
    SRMux I__1160 (
            .O(N__5850),
            .I(N__5664));
    SRMux I__1159 (
            .O(N__5849),
            .I(N__5664));
    SRMux I__1158 (
            .O(N__5848),
            .I(N__5664));
    SRMux I__1157 (
            .O(N__5847),
            .I(N__5664));
    SRMux I__1156 (
            .O(N__5846),
            .I(N__5664));
    SRMux I__1155 (
            .O(N__5845),
            .I(N__5664));
    SRMux I__1154 (
            .O(N__5844),
            .I(N__5664));
    SRMux I__1153 (
            .O(N__5843),
            .I(N__5664));
    SRMux I__1152 (
            .O(N__5842),
            .I(N__5664));
    SRMux I__1151 (
            .O(N__5841),
            .I(N__5664));
    SRMux I__1150 (
            .O(N__5840),
            .I(N__5664));
    SRMux I__1149 (
            .O(N__5839),
            .I(N__5664));
    SRMux I__1148 (
            .O(N__5838),
            .I(N__5664));
    SRMux I__1147 (
            .O(N__5837),
            .I(N__5664));
    SRMux I__1146 (
            .O(N__5836),
            .I(N__5664));
    SRMux I__1145 (
            .O(N__5835),
            .I(N__5664));
    SRMux I__1144 (
            .O(N__5834),
            .I(N__5664));
    SRMux I__1143 (
            .O(N__5833),
            .I(N__5664));
    SRMux I__1142 (
            .O(N__5832),
            .I(N__5664));
    SRMux I__1141 (
            .O(N__5831),
            .I(N__5664));
    SRMux I__1140 (
            .O(N__5830),
            .I(N__5664));
    SRMux I__1139 (
            .O(N__5829),
            .I(N__5664));
    SRMux I__1138 (
            .O(N__5828),
            .I(N__5664));
    SRMux I__1137 (
            .O(N__5827),
            .I(N__5664));
    SRMux I__1136 (
            .O(N__5826),
            .I(N__5664));
    SRMux I__1135 (
            .O(N__5825),
            .I(N__5664));
    SRMux I__1134 (
            .O(N__5824),
            .I(N__5664));
    SRMux I__1133 (
            .O(N__5823),
            .I(N__5664));
    SRMux I__1132 (
            .O(N__5822),
            .I(N__5664));
    SRMux I__1131 (
            .O(N__5821),
            .I(N__5664));
    SRMux I__1130 (
            .O(N__5820),
            .I(N__5664));
    SRMux I__1129 (
            .O(N__5819),
            .I(N__5664));
    SRMux I__1128 (
            .O(N__5818),
            .I(N__5664));
    SRMux I__1127 (
            .O(N__5817),
            .I(N__5664));
    SRMux I__1126 (
            .O(N__5816),
            .I(N__5664));
    SRMux I__1125 (
            .O(N__5815),
            .I(N__5664));
    SRMux I__1124 (
            .O(N__5814),
            .I(N__5664));
    SRMux I__1123 (
            .O(N__5813),
            .I(N__5664));
    SRMux I__1122 (
            .O(N__5812),
            .I(N__5664));
    SRMux I__1121 (
            .O(N__5811),
            .I(N__5664));
    SRMux I__1120 (
            .O(N__5810),
            .I(N__5664));
    SRMux I__1119 (
            .O(N__5809),
            .I(N__5664));
    SRMux I__1118 (
            .O(N__5808),
            .I(N__5664));
    SRMux I__1117 (
            .O(N__5807),
            .I(N__5664));
    SRMux I__1116 (
            .O(N__5806),
            .I(N__5664));
    SRMux I__1115 (
            .O(N__5805),
            .I(N__5664));
    SRMux I__1114 (
            .O(N__5804),
            .I(N__5664));
    SRMux I__1113 (
            .O(N__5803),
            .I(N__5664));
    SRMux I__1112 (
            .O(N__5802),
            .I(N__5664));
    SRMux I__1111 (
            .O(N__5801),
            .I(N__5664));
    GlobalMux I__1110 (
            .O(N__5664),
            .I(N__5661));
    gio2CtrlBuf I__1109 (
            .O(N__5661),
            .I(RST_N_c_i_g));
    InMux I__1108 (
            .O(N__5658),
            .I(N__5655));
    LocalMux I__1107 (
            .O(N__5655),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_61 ));
    InMux I__1106 (
            .O(N__5652),
            .I(N__5649));
    LocalMux I__1105 (
            .O(N__5649),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_62 ));
    InMux I__1104 (
            .O(N__5646),
            .I(N__5643));
    LocalMux I__1103 (
            .O(N__5643),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_30 ));
    InMux I__1102 (
            .O(N__5640),
            .I(N__5637));
    LocalMux I__1101 (
            .O(N__5637),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_34 ));
    InMux I__1100 (
            .O(N__5634),
            .I(N__5631));
    LocalMux I__1099 (
            .O(N__5631),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_31 ));
    InMux I__1098 (
            .O(N__5628),
            .I(N__5625));
    LocalMux I__1097 (
            .O(N__5625),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_32 ));
    InMux I__1096 (
            .O(N__5622),
            .I(N__5619));
    LocalMux I__1095 (
            .O(N__5619),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_33 ));
    InMux I__1094 (
            .O(N__5616),
            .I(N__5613));
    LocalMux I__1093 (
            .O(N__5613),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_26 ));
    InMux I__1092 (
            .O(N__5610),
            .I(N__5607));
    LocalMux I__1091 (
            .O(N__5607),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_24 ));
    InMux I__1090 (
            .O(N__5604),
            .I(N__5601));
    LocalMux I__1089 (
            .O(N__5601),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_25 ));
    InMux I__1088 (
            .O(N__5598),
            .I(N__5595));
    LocalMux I__1087 (
            .O(N__5595),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_23 ));
    InMux I__1086 (
            .O(N__5592),
            .I(N__5589));
    LocalMux I__1085 (
            .O(N__5589),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_49 ));
    InMux I__1084 (
            .O(N__5586),
            .I(N__5583));
    LocalMux I__1083 (
            .O(N__5583),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_52 ));
    InMux I__1082 (
            .O(N__5580),
            .I(N__5577));
    LocalMux I__1081 (
            .O(N__5577),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_50 ));
    InMux I__1080 (
            .O(N__5574),
            .I(N__5571));
    LocalMux I__1079 (
            .O(N__5571),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_51 ));
    InMux I__1078 (
            .O(N__5568),
            .I(N__5565));
    LocalMux I__1077 (
            .O(N__5565),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_64 ));
    InMux I__1076 (
            .O(N__5562),
            .I(N__5559));
    LocalMux I__1075 (
            .O(N__5559),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_63 ));
    InMux I__1074 (
            .O(N__5556),
            .I(N__5553));
    LocalMux I__1073 (
            .O(N__5553),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_53 ));
    InMux I__1072 (
            .O(N__5550),
            .I(N__5547));
    LocalMux I__1071 (
            .O(N__5547),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_36 ));
    InMux I__1070 (
            .O(N__5544),
            .I(N__5541));
    LocalMux I__1069 (
            .O(N__5541),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_35 ));
    InMux I__1068 (
            .O(N__5538),
            .I(N__5535));
    LocalMux I__1067 (
            .O(N__5535),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_37 ));
    InMux I__1066 (
            .O(N__5532),
            .I(N__5529));
    LocalMux I__1065 (
            .O(N__5529),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_38 ));
    InMux I__1064 (
            .O(N__5526),
            .I(N__5523));
    LocalMux I__1063 (
            .O(N__5523),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_39 ));
    InMux I__1062 (
            .O(N__5520),
            .I(N__5517));
    LocalMux I__1061 (
            .O(N__5517),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_46 ));
    InMux I__1060 (
            .O(N__5514),
            .I(N__5511));
    LocalMux I__1059 (
            .O(N__5511),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_47 ));
    InMux I__1058 (
            .O(N__5508),
            .I(N__5505));
    LocalMux I__1057 (
            .O(N__5505),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_22 ));
    InMux I__1056 (
            .O(N__5502),
            .I(N__5499));
    LocalMux I__1055 (
            .O(N__5499),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_48 ));
    InMux I__1054 (
            .O(N__5496),
            .I(N__5493));
    LocalMux I__1053 (
            .O(N__5493),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_19 ));
    InMux I__1052 (
            .O(N__5490),
            .I(N__5487));
    LocalMux I__1051 (
            .O(N__5487),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_20 ));
    InMux I__1050 (
            .O(N__5484),
            .I(N__5481));
    LocalMux I__1049 (
            .O(N__5481),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_41 ));
    InMux I__1048 (
            .O(N__5478),
            .I(N__5475));
    LocalMux I__1047 (
            .O(N__5475),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_40 ));
    InMux I__1046 (
            .O(N__5472),
            .I(N__5469));
    LocalMux I__1045 (
            .O(N__5469),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_42 ));
    InMux I__1044 (
            .O(N__5466),
            .I(N__5463));
    LocalMux I__1043 (
            .O(N__5463),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_43 ));
    InMux I__1042 (
            .O(N__5460),
            .I(N__5457));
    LocalMux I__1041 (
            .O(N__5457),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_44 ));
    InMux I__1040 (
            .O(N__5454),
            .I(N__5451));
    LocalMux I__1039 (
            .O(N__5451),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_45 ));
    InMux I__1038 (
            .O(N__5448),
            .I(N__5445));
    LocalMux I__1037 (
            .O(N__5445),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_21 ));
    InMux I__1036 (
            .O(N__5442),
            .I(N__5439));
    LocalMux I__1035 (
            .O(N__5439),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_65 ));
    InMux I__1034 (
            .O(N__5436),
            .I(N__5433));
    LocalMux I__1033 (
            .O(N__5433),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_18 ));
    InMux I__1032 (
            .O(N__5430),
            .I(N__5427));
    LocalMux I__1031 (
            .O(N__5427),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_71 ));
    InMux I__1030 (
            .O(N__5424),
            .I(N__5421));
    LocalMux I__1029 (
            .O(N__5421),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_72 ));
    InMux I__1028 (
            .O(N__5418),
            .I(N__5415));
    LocalMux I__1027 (
            .O(N__5415),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_70 ));
    InMux I__1026 (
            .O(N__5412),
            .I(N__5409));
    LocalMux I__1025 (
            .O(N__5409),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_68 ));
    InMux I__1024 (
            .O(N__5406),
            .I(N__5403));
    LocalMux I__1023 (
            .O(N__5403),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_69 ));
    InMux I__1022 (
            .O(N__5400),
            .I(N__5397));
    LocalMux I__1021 (
            .O(N__5397),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_67 ));
    InMux I__1020 (
            .O(N__5394),
            .I(N__5391));
    LocalMux I__1019 (
            .O(N__5391),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_66 ));
    InMux I__1018 (
            .O(N__5388),
            .I(N__5385));
    LocalMux I__1017 (
            .O(N__5385),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_77 ));
    InMux I__1016 (
            .O(N__5382),
            .I(N__5379));
    LocalMux I__1015 (
            .O(N__5379),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_78 ));
    InMux I__1014 (
            .O(N__5376),
            .I(N__5373));
    LocalMux I__1013 (
            .O(N__5373),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_14 ));
    InMux I__1012 (
            .O(N__5370),
            .I(N__5367));
    LocalMux I__1011 (
            .O(N__5367),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_75 ));
    InMux I__1010 (
            .O(N__5364),
            .I(N__5361));
    LocalMux I__1009 (
            .O(N__5361),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_76 ));
    InMux I__1008 (
            .O(N__5358),
            .I(N__5355));
    LocalMux I__1007 (
            .O(N__5355),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_74 ));
    InMux I__1006 (
            .O(N__5352),
            .I(N__5349));
    LocalMux I__1005 (
            .O(N__5349),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_15 ));
    InMux I__1004 (
            .O(N__5346),
            .I(N__5343));
    LocalMux I__1003 (
            .O(N__5343),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_16 ));
    InMux I__1002 (
            .O(N__5340),
            .I(N__5337));
    LocalMux I__1001 (
            .O(N__5337),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_73 ));
    InMux I__1000 (
            .O(N__5334),
            .I(N__5331));
    LocalMux I__999 (
            .O(N__5331),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_17 ));
    InMux I__998 (
            .O(N__5328),
            .I(N__5325));
    LocalMux I__997 (
            .O(N__5325),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_10 ));
    InMux I__996 (
            .O(N__5322),
            .I(N__5319));
    LocalMux I__995 (
            .O(N__5319),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_11 ));
    InMux I__994 (
            .O(N__5316),
            .I(N__5313));
    LocalMux I__993 (
            .O(N__5313),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_83 ));
    InMux I__992 (
            .O(N__5310),
            .I(N__5307));
    LocalMux I__991 (
            .O(N__5307),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_12 ));
    InMux I__990 (
            .O(N__5304),
            .I(N__5301));
    LocalMux I__989 (
            .O(N__5301),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_81 ));
    InMux I__988 (
            .O(N__5298),
            .I(N__5295));
    LocalMux I__987 (
            .O(N__5295),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_82 ));
    InMux I__986 (
            .O(N__5292),
            .I(N__5289));
    LocalMux I__985 (
            .O(N__5289),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_13 ));
    InMux I__984 (
            .O(N__5286),
            .I(N__5283));
    LocalMux I__983 (
            .O(N__5283),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_80 ));
    InMux I__982 (
            .O(N__5280),
            .I(N__5277));
    LocalMux I__981 (
            .O(N__5277),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_79 ));
    InMux I__980 (
            .O(N__5274),
            .I(N__5271));
    LocalMux I__979 (
            .O(N__5271),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_4 ));
    InMux I__978 (
            .O(N__5268),
            .I(N__5265));
    LocalMux I__977 (
            .O(N__5265),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_5 ));
    InMux I__976 (
            .O(N__5262),
            .I(N__5259));
    LocalMux I__975 (
            .O(N__5259),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_86 ));
    InMux I__974 (
            .O(N__5256),
            .I(N__5253));
    LocalMux I__973 (
            .O(N__5253),
            .I(N__5250));
    Odrv4 I__972 (
            .O(N__5250),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_6 ));
    InMux I__971 (
            .O(N__5247),
            .I(N__5244));
    LocalMux I__970 (
            .O(N__5244),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_7 ));
    InMux I__969 (
            .O(N__5241),
            .I(N__5238));
    LocalMux I__968 (
            .O(N__5238),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_8 ));
    InMux I__967 (
            .O(N__5235),
            .I(N__5232));
    LocalMux I__966 (
            .O(N__5232),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_84 ));
    InMux I__965 (
            .O(N__5229),
            .I(N__5226));
    LocalMux I__964 (
            .O(N__5226),
            .I(N__5223));
    Odrv4 I__963 (
            .O(N__5223),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_85 ));
    InMux I__962 (
            .O(N__5220),
            .I(N__5217));
    LocalMux I__961 (
            .O(N__5217),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_9 ));
    InMux I__960 (
            .O(N__5214),
            .I(N__5211));
    LocalMux I__959 (
            .O(N__5211),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_2 ));
    InMux I__958 (
            .O(N__5208),
            .I(N__5205));
    LocalMux I__957 (
            .O(N__5205),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_3 ));
    InMux I__956 (
            .O(N__5202),
            .I(N__5199));
    LocalMux I__955 (
            .O(N__5199),
            .I(N__5196));
    Odrv12 I__954 (
            .O(N__5196),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_87 ));
    InMux I__953 (
            .O(N__5193),
            .I(N__5190));
    LocalMux I__952 (
            .O(N__5190),
            .I(\config_register_latched_dec_inst1.DYNSRZ0Z_9 ));
    InMux I__951 (
            .O(N__5187),
            .I(N__5184));
    LocalMux I__950 (
            .O(N__5184),
            .I(\config_register_latched_dec_inst1.DYNSRZ0Z_6 ));
    InMux I__949 (
            .O(N__5181),
            .I(N__5178));
    LocalMux I__948 (
            .O(N__5178),
            .I(\config_register_latched_dec_inst1.DYNSRZ0Z_7 ));
    InMux I__947 (
            .O(N__5175),
            .I(N__5172));
    LocalMux I__946 (
            .O(N__5172),
            .I(\config_register_latched_dec_inst1.DYNSRZ0Z_8 ));
    InMux I__945 (
            .O(N__5169),
            .I(N__5166));
    LocalMux I__944 (
            .O(N__5166),
            .I(\config_register_latched_dec_inst1.DYNSRZ0Z_4 ));
    InMux I__943 (
            .O(N__5163),
            .I(N__5160));
    LocalMux I__942 (
            .O(N__5160),
            .I(\config_register_latched_dec_inst1.DYNSRZ0Z_5 ));
    CEMux I__941 (
            .O(N__5157),
            .I(N__5154));
    LocalMux I__940 (
            .O(N__5154),
            .I(N__5149));
    CEMux I__939 (
            .O(N__5153),
            .I(N__5146));
    CEMux I__938 (
            .O(N__5152),
            .I(N__5142));
    Span4Mux_h I__937 (
            .O(N__5149),
            .I(N__5137));
    LocalMux I__936 (
            .O(N__5146),
            .I(N__5137));
    CEMux I__935 (
            .O(N__5145),
            .I(N__5134));
    LocalMux I__934 (
            .O(N__5142),
            .I(N__5131));
    Span4Mux_v I__933 (
            .O(N__5137),
            .I(N__5126));
    LocalMux I__932 (
            .O(N__5134),
            .I(N__5126));
    Span4Mux_h I__931 (
            .O(N__5131),
            .I(N__5123));
    Span4Mux_v I__930 (
            .O(N__5126),
            .I(N__5120));
    Odrv4 I__929 (
            .O(N__5123),
            .I(\config_register_latched_dec_inst1.DYNSR_cnv_nsZ0Z_0 ));
    Odrv4 I__928 (
            .O(N__5120),
            .I(\config_register_latched_dec_inst1.DYNSR_cnv_nsZ0Z_0 ));
    CascadeMux I__927 (
            .O(N__5115),
            .I(N__5109));
    InMux I__926 (
            .O(N__5114),
            .I(N__5106));
    InMux I__925 (
            .O(N__5113),
            .I(N__5099));
    InMux I__924 (
            .O(N__5112),
            .I(N__5099));
    InMux I__923 (
            .O(N__5109),
            .I(N__5099));
    LocalMux I__922 (
            .O(N__5106),
            .I(N__5094));
    LocalMux I__921 (
            .O(N__5099),
            .I(N__5094));
    Span4Mux_v I__920 (
            .O(N__5094),
            .I(N__5090));
    InMux I__919 (
            .O(N__5093),
            .I(N__5087));
    Span4Mux_h I__918 (
            .O(N__5090),
            .I(N__5084));
    LocalMux I__917 (
            .O(N__5087),
            .I(N__5081));
    Odrv4 I__916 (
            .O(N__5084),
            .I(CLK_uC_c));
    Odrv12 I__915 (
            .O(N__5081),
            .I(CLK_uC_c));
    CascadeMux I__914 (
            .O(N__5076),
            .I(N__5070));
    InMux I__913 (
            .O(N__5075),
            .I(N__5063));
    InMux I__912 (
            .O(N__5074),
            .I(N__5063));
    InMux I__911 (
            .O(N__5073),
            .I(N__5063));
    InMux I__910 (
            .O(N__5070),
            .I(N__5060));
    LocalMux I__909 (
            .O(N__5063),
            .I(fsm_ctrl_inst1_SCLK_i));
    LocalMux I__908 (
            .O(N__5060),
            .I(fsm_ctrl_inst1_SCLK_i));
    InMux I__907 (
            .O(N__5055),
            .I(N__5040));
    InMux I__906 (
            .O(N__5054),
            .I(N__5040));
    InMux I__905 (
            .O(N__5053),
            .I(N__5025));
    InMux I__904 (
            .O(N__5052),
            .I(N__5025));
    InMux I__903 (
            .O(N__5051),
            .I(N__5025));
    InMux I__902 (
            .O(N__5050),
            .I(N__5025));
    InMux I__901 (
            .O(N__5049),
            .I(N__5025));
    InMux I__900 (
            .O(N__5048),
            .I(N__5019));
    InMux I__899 (
            .O(N__5047),
            .I(N__5012));
    InMux I__898 (
            .O(N__5046),
            .I(N__5012));
    InMux I__897 (
            .O(N__5045),
            .I(N__5012));
    LocalMux I__896 (
            .O(N__5040),
            .I(N__4980));
    InMux I__895 (
            .O(N__5039),
            .I(N__4973));
    InMux I__894 (
            .O(N__5038),
            .I(N__4973));
    InMux I__893 (
            .O(N__5037),
            .I(N__4973));
    InMux I__892 (
            .O(N__5036),
            .I(N__4957));
    LocalMux I__891 (
            .O(N__5025),
            .I(N__4939));
    InMux I__890 (
            .O(N__5024),
            .I(N__4932));
    InMux I__889 (
            .O(N__5023),
            .I(N__4932));
    InMux I__888 (
            .O(N__5022),
            .I(N__4932));
    LocalMux I__887 (
            .O(N__5019),
            .I(N__4927));
    LocalMux I__886 (
            .O(N__5012),
            .I(N__4927));
    InMux I__885 (
            .O(N__5011),
            .I(N__4922));
    InMux I__884 (
            .O(N__5010),
            .I(N__4922));
    InMux I__883 (
            .O(N__5009),
            .I(N__4911));
    InMux I__882 (
            .O(N__5008),
            .I(N__4911));
    InMux I__881 (
            .O(N__5007),
            .I(N__4911));
    InMux I__880 (
            .O(N__5006),
            .I(N__4911));
    InMux I__879 (
            .O(N__5005),
            .I(N__4911));
    InMux I__878 (
            .O(N__5004),
            .I(N__4900));
    InMux I__877 (
            .O(N__5003),
            .I(N__4900));
    InMux I__876 (
            .O(N__5002),
            .I(N__4900));
    InMux I__875 (
            .O(N__5001),
            .I(N__4900));
    InMux I__874 (
            .O(N__5000),
            .I(N__4900));
    InMux I__873 (
            .O(N__4999),
            .I(N__4885));
    InMux I__872 (
            .O(N__4998),
            .I(N__4885));
    InMux I__871 (
            .O(N__4997),
            .I(N__4885));
    InMux I__870 (
            .O(N__4996),
            .I(N__4885));
    InMux I__869 (
            .O(N__4995),
            .I(N__4885));
    InMux I__868 (
            .O(N__4994),
            .I(N__4885));
    InMux I__867 (
            .O(N__4993),
            .I(N__4885));
    InMux I__866 (
            .O(N__4992),
            .I(N__4868));
    InMux I__865 (
            .O(N__4991),
            .I(N__4868));
    InMux I__864 (
            .O(N__4990),
            .I(N__4868));
    InMux I__863 (
            .O(N__4989),
            .I(N__4868));
    InMux I__862 (
            .O(N__4988),
            .I(N__4868));
    InMux I__861 (
            .O(N__4987),
            .I(N__4868));
    InMux I__860 (
            .O(N__4986),
            .I(N__4868));
    InMux I__859 (
            .O(N__4985),
            .I(N__4868));
    InMux I__858 (
            .O(N__4984),
            .I(N__4847));
    InMux I__857 (
            .O(N__4983),
            .I(N__4847));
    Span4Mux_s2_h I__856 (
            .O(N__4980),
            .I(N__4842));
    LocalMux I__855 (
            .O(N__4973),
            .I(N__4842));
    InMux I__854 (
            .O(N__4972),
            .I(N__4839));
    InMux I__853 (
            .O(N__4971),
            .I(N__4828));
    InMux I__852 (
            .O(N__4970),
            .I(N__4828));
    InMux I__851 (
            .O(N__4969),
            .I(N__4828));
    InMux I__850 (
            .O(N__4968),
            .I(N__4828));
    InMux I__849 (
            .O(N__4967),
            .I(N__4828));
    InMux I__848 (
            .O(N__4966),
            .I(N__4823));
    InMux I__847 (
            .O(N__4965),
            .I(N__4823));
    InMux I__846 (
            .O(N__4964),
            .I(N__4814));
    InMux I__845 (
            .O(N__4963),
            .I(N__4814));
    InMux I__844 (
            .O(N__4962),
            .I(N__4814));
    InMux I__843 (
            .O(N__4961),
            .I(N__4814));
    CascadeMux I__842 (
            .O(N__4960),
            .I(N__4811));
    LocalMux I__841 (
            .O(N__4957),
            .I(N__4803));
    InMux I__840 (
            .O(N__4956),
            .I(N__4788));
    InMux I__839 (
            .O(N__4955),
            .I(N__4788));
    InMux I__838 (
            .O(N__4954),
            .I(N__4788));
    InMux I__837 (
            .O(N__4953),
            .I(N__4788));
    InMux I__836 (
            .O(N__4952),
            .I(N__4788));
    InMux I__835 (
            .O(N__4951),
            .I(N__4788));
    InMux I__834 (
            .O(N__4950),
            .I(N__4788));
    InMux I__833 (
            .O(N__4949),
            .I(N__4771));
    InMux I__832 (
            .O(N__4948),
            .I(N__4771));
    InMux I__831 (
            .O(N__4947),
            .I(N__4771));
    InMux I__830 (
            .O(N__4946),
            .I(N__4771));
    InMux I__829 (
            .O(N__4945),
            .I(N__4771));
    InMux I__828 (
            .O(N__4944),
            .I(N__4771));
    InMux I__827 (
            .O(N__4943),
            .I(N__4771));
    InMux I__826 (
            .O(N__4942),
            .I(N__4771));
    Span4Mux_v I__825 (
            .O(N__4939),
            .I(N__4756));
    LocalMux I__824 (
            .O(N__4932),
            .I(N__4756));
    Span4Mux_h I__823 (
            .O(N__4927),
            .I(N__4756));
    LocalMux I__822 (
            .O(N__4922),
            .I(N__4756));
    LocalMux I__821 (
            .O(N__4911),
            .I(N__4756));
    LocalMux I__820 (
            .O(N__4900),
            .I(N__4756));
    LocalMux I__819 (
            .O(N__4885),
            .I(N__4756));
    LocalMux I__818 (
            .O(N__4868),
            .I(N__4753));
    InMux I__817 (
            .O(N__4867),
            .I(N__4738));
    InMux I__816 (
            .O(N__4866),
            .I(N__4738));
    InMux I__815 (
            .O(N__4865),
            .I(N__4738));
    InMux I__814 (
            .O(N__4864),
            .I(N__4738));
    InMux I__813 (
            .O(N__4863),
            .I(N__4738));
    InMux I__812 (
            .O(N__4862),
            .I(N__4738));
    InMux I__811 (
            .O(N__4861),
            .I(N__4738));
    InMux I__810 (
            .O(N__4860),
            .I(N__4721));
    InMux I__809 (
            .O(N__4859),
            .I(N__4721));
    InMux I__808 (
            .O(N__4858),
            .I(N__4721));
    InMux I__807 (
            .O(N__4857),
            .I(N__4721));
    InMux I__806 (
            .O(N__4856),
            .I(N__4721));
    InMux I__805 (
            .O(N__4855),
            .I(N__4721));
    InMux I__804 (
            .O(N__4854),
            .I(N__4721));
    InMux I__803 (
            .O(N__4853),
            .I(N__4721));
    InMux I__802 (
            .O(N__4852),
            .I(N__4718));
    LocalMux I__801 (
            .O(N__4847),
            .I(N__4707));
    Span4Mux_h I__800 (
            .O(N__4842),
            .I(N__4707));
    LocalMux I__799 (
            .O(N__4839),
            .I(N__4707));
    LocalMux I__798 (
            .O(N__4828),
            .I(N__4707));
    LocalMux I__797 (
            .O(N__4823),
            .I(N__4707));
    LocalMux I__796 (
            .O(N__4814),
            .I(N__4704));
    InMux I__795 (
            .O(N__4811),
            .I(N__4701));
    CascadeMux I__794 (
            .O(N__4810),
            .I(N__4698));
    CascadeMux I__793 (
            .O(N__4809),
            .I(N__4695));
    CascadeMux I__792 (
            .O(N__4808),
            .I(N__4691));
    InMux I__791 (
            .O(N__4807),
            .I(N__4684));
    InMux I__790 (
            .O(N__4806),
            .I(N__4681));
    Span12Mux_s4_h I__789 (
            .O(N__4803),
            .I(N__4674));
    LocalMux I__788 (
            .O(N__4788),
            .I(N__4674));
    LocalMux I__787 (
            .O(N__4771),
            .I(N__4674));
    Span4Mux_v I__786 (
            .O(N__4756),
            .I(N__4665));
    Span4Mux_h I__785 (
            .O(N__4753),
            .I(N__4665));
    LocalMux I__784 (
            .O(N__4738),
            .I(N__4665));
    LocalMux I__783 (
            .O(N__4721),
            .I(N__4665));
    LocalMux I__782 (
            .O(N__4718),
            .I(N__4656));
    Span4Mux_v I__781 (
            .O(N__4707),
            .I(N__4656));
    Span4Mux_s2_h I__780 (
            .O(N__4704),
            .I(N__4656));
    LocalMux I__779 (
            .O(N__4701),
            .I(N__4656));
    InMux I__778 (
            .O(N__4698),
            .I(N__4651));
    InMux I__777 (
            .O(N__4695),
            .I(N__4651));
    InMux I__776 (
            .O(N__4694),
            .I(N__4648));
    InMux I__775 (
            .O(N__4691),
            .I(N__4643));
    InMux I__774 (
            .O(N__4690),
            .I(N__4643));
    InMux I__773 (
            .O(N__4689),
            .I(N__4636));
    InMux I__772 (
            .O(N__4688),
            .I(N__4636));
    InMux I__771 (
            .O(N__4687),
            .I(N__4636));
    LocalMux I__770 (
            .O(N__4684),
            .I(fsm_ctrl_inst1_current_state_1));
    LocalMux I__769 (
            .O(N__4681),
            .I(fsm_ctrl_inst1_current_state_1));
    Odrv12 I__768 (
            .O(N__4674),
            .I(fsm_ctrl_inst1_current_state_1));
    Odrv4 I__767 (
            .O(N__4665),
            .I(fsm_ctrl_inst1_current_state_1));
    Odrv4 I__766 (
            .O(N__4656),
            .I(fsm_ctrl_inst1_current_state_1));
    LocalMux I__765 (
            .O(N__4651),
            .I(fsm_ctrl_inst1_current_state_1));
    LocalMux I__764 (
            .O(N__4648),
            .I(fsm_ctrl_inst1_current_state_1));
    LocalMux I__763 (
            .O(N__4643),
            .I(fsm_ctrl_inst1_current_state_1));
    LocalMux I__762 (
            .O(N__4636),
            .I(fsm_ctrl_inst1_current_state_1));
    CascadeMux I__761 (
            .O(N__4617),
            .I(\config_register_latched_dec_inst1.STATSR_cnv_x1Z0Z_0_cascade_ ));
    InMux I__760 (
            .O(N__4614),
            .I(N__4611));
    LocalMux I__759 (
            .O(N__4611),
            .I(\config_register_latched_dec_inst1.STATSR_cnv_x0Z0Z_0 ));
    IoInMux I__758 (
            .O(N__4608),
            .I(N__4605));
    LocalMux I__757 (
            .O(N__4605),
            .I(N__4602));
    Span12Mux_s11_v I__756 (
            .O(N__4602),
            .I(N__4599));
    Odrv12 I__755 (
            .O(N__4599),
            .I(STATSR_cnv_ns_0));
    InMux I__754 (
            .O(N__4596),
            .I(N__4585));
    InMux I__753 (
            .O(N__4595),
            .I(N__4570));
    InMux I__752 (
            .O(N__4594),
            .I(N__4570));
    InMux I__751 (
            .O(N__4593),
            .I(N__4570));
    InMux I__750 (
            .O(N__4592),
            .I(N__4570));
    InMux I__749 (
            .O(N__4591),
            .I(N__4570));
    InMux I__748 (
            .O(N__4590),
            .I(N__4570));
    InMux I__747 (
            .O(N__4589),
            .I(N__4560));
    InMux I__746 (
            .O(N__4588),
            .I(N__4560));
    LocalMux I__745 (
            .O(N__4585),
            .I(N__4557));
    InMux I__744 (
            .O(N__4584),
            .I(N__4536));
    InMux I__743 (
            .O(N__4583),
            .I(N__4536));
    LocalMux I__742 (
            .O(N__4570),
            .I(N__4533));
    InMux I__741 (
            .O(N__4569),
            .I(N__4522));
    InMux I__740 (
            .O(N__4568),
            .I(N__4522));
    InMux I__739 (
            .O(N__4567),
            .I(N__4522));
    InMux I__738 (
            .O(N__4566),
            .I(N__4522));
    InMux I__737 (
            .O(N__4565),
            .I(N__4522));
    LocalMux I__736 (
            .O(N__4560),
            .I(N__4517));
    Span4Mux_s2_h I__735 (
            .O(N__4557),
            .I(N__4517));
    InMux I__734 (
            .O(N__4556),
            .I(N__4510));
    InMux I__733 (
            .O(N__4555),
            .I(N__4510));
    InMux I__732 (
            .O(N__4554),
            .I(N__4510));
    InMux I__731 (
            .O(N__4553),
            .I(N__4504));
    InMux I__730 (
            .O(N__4552),
            .I(N__4487));
    InMux I__729 (
            .O(N__4551),
            .I(N__4487));
    InMux I__728 (
            .O(N__4550),
            .I(N__4487));
    InMux I__727 (
            .O(N__4549),
            .I(N__4487));
    InMux I__726 (
            .O(N__4548),
            .I(N__4487));
    InMux I__725 (
            .O(N__4547),
            .I(N__4487));
    InMux I__724 (
            .O(N__4546),
            .I(N__4487));
    InMux I__723 (
            .O(N__4545),
            .I(N__4487));
    InMux I__722 (
            .O(N__4544),
            .I(N__4482));
    InMux I__721 (
            .O(N__4543),
            .I(N__4482));
    InMux I__720 (
            .O(N__4542),
            .I(N__4477));
    InMux I__719 (
            .O(N__4541),
            .I(N__4477));
    LocalMux I__718 (
            .O(N__4536),
            .I(N__4466));
    Span4Mux_v I__717 (
            .O(N__4533),
            .I(N__4466));
    LocalMux I__716 (
            .O(N__4522),
            .I(N__4466));
    Span4Mux_v I__715 (
            .O(N__4517),
            .I(N__4466));
    LocalMux I__714 (
            .O(N__4510),
            .I(N__4466));
    InMux I__713 (
            .O(N__4509),
            .I(N__4459));
    InMux I__712 (
            .O(N__4508),
            .I(N__4459));
    InMux I__711 (
            .O(N__4507),
            .I(N__4459));
    LocalMux I__710 (
            .O(N__4504),
            .I(fsm_ctrl_inst1_current_state_0));
    LocalMux I__709 (
            .O(N__4487),
            .I(fsm_ctrl_inst1_current_state_0));
    LocalMux I__708 (
            .O(N__4482),
            .I(fsm_ctrl_inst1_current_state_0));
    LocalMux I__707 (
            .O(N__4477),
            .I(fsm_ctrl_inst1_current_state_0));
    Odrv4 I__706 (
            .O(N__4466),
            .I(fsm_ctrl_inst1_current_state_0));
    LocalMux I__705 (
            .O(N__4459),
            .I(fsm_ctrl_inst1_current_state_0));
    InMux I__704 (
            .O(N__4446),
            .I(N__4443));
    LocalMux I__703 (
            .O(N__4443),
            .I(N__4436));
    InMux I__702 (
            .O(N__4442),
            .I(N__4429));
    InMux I__701 (
            .O(N__4441),
            .I(N__4429));
    InMux I__700 (
            .O(N__4440),
            .I(N__4429));
    InMux I__699 (
            .O(N__4439),
            .I(N__4426));
    Odrv4 I__698 (
            .O(N__4436),
            .I(SEL_REG));
    LocalMux I__697 (
            .O(N__4429),
            .I(SEL_REG));
    LocalMux I__696 (
            .O(N__4426),
            .I(SEL_REG));
    InMux I__695 (
            .O(N__4419),
            .I(N__4415));
    InMux I__694 (
            .O(N__4418),
            .I(N__4412));
    LocalMux I__693 (
            .O(N__4415),
            .I(N__4409));
    LocalMux I__692 (
            .O(N__4412),
            .I(MOSI));
    Odrv4 I__691 (
            .O(N__4409),
            .I(MOSI));
    InMux I__690 (
            .O(N__4404),
            .I(N__4401));
    LocalMux I__689 (
            .O(N__4401),
            .I(\config_register_latched_dec_inst1.DYNSRZ0Z_0 ));
    InMux I__688 (
            .O(N__4398),
            .I(N__4395));
    LocalMux I__687 (
            .O(N__4395),
            .I(\config_register_latched_dec_inst1.DYNSRZ0Z_1 ));
    InMux I__686 (
            .O(N__4392),
            .I(N__4389));
    LocalMux I__685 (
            .O(N__4389),
            .I(\config_register_latched_dec_inst1.DYNSRZ0Z_2 ));
    InMux I__684 (
            .O(N__4386),
            .I(N__4383));
    LocalMux I__683 (
            .O(N__4383),
            .I(\config_register_latched_dec_inst1.DYNSRZ0Z_3 ));
    InMux I__682 (
            .O(N__4380),
            .I(N__4377));
    LocalMux I__681 (
            .O(N__4377),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_1 ));
    InMux I__680 (
            .O(N__4374),
            .I(N__4371));
    LocalMux I__679 (
            .O(N__4371),
            .I(\config_register_latched_dec_inst1.DYNSRZ0Z_14 ));
    InMux I__678 (
            .O(N__4368),
            .I(N__4365));
    LocalMux I__677 (
            .O(N__4365),
            .I(\config_register_latched_dec_inst1.DYNSRZ0Z_15 ));
    InMux I__676 (
            .O(N__4362),
            .I(N__4359));
    LocalMux I__675 (
            .O(N__4359),
            .I(\config_register_latched_dec_inst1.DYNSRZ0Z_12 ));
    InMux I__674 (
            .O(N__4356),
            .I(N__4353));
    LocalMux I__673 (
            .O(N__4353),
            .I(\config_register_latched_dec_inst1.DYNSRZ0Z_13 ));
    InMux I__672 (
            .O(N__4350),
            .I(N__4347));
    LocalMux I__671 (
            .O(N__4347),
            .I(\config_register_latched_dec_inst1.DYNSRZ0Z_10 ));
    InMux I__670 (
            .O(N__4344),
            .I(N__4341));
    LocalMux I__669 (
            .O(N__4341),
            .I(\config_register_latched_dec_inst1.DYNSRZ0Z_11 ));
    CascadeMux I__668 (
            .O(N__4338),
            .I(\config_register_latched_dec_inst1.DYNSR_cnv_x0Z0Z_0_cascade_ ));
    InMux I__667 (
            .O(N__4335),
            .I(N__4332));
    LocalMux I__666 (
            .O(N__4332),
            .I(\config_register_latched_dec_inst1.DYNSR_cnv_x1Z0Z_0 ));
    InMux I__665 (
            .O(N__4329),
            .I(N__4317));
    InMux I__664 (
            .O(N__4328),
            .I(N__4317));
    InMux I__663 (
            .O(N__4327),
            .I(N__4317));
    InMux I__662 (
            .O(N__4326),
            .I(N__4317));
    LocalMux I__661 (
            .O(N__4317),
            .I(\fsm_ctrl_inst1.counter_dinZ0Z_2 ));
    CascadeMux I__660 (
            .O(N__4314),
            .I(N__4309));
    CascadeMux I__659 (
            .O(N__4313),
            .I(N__4306));
    CascadeMux I__658 (
            .O(N__4312),
            .I(N__4303));
    InMux I__657 (
            .O(N__4309),
            .I(N__4296));
    InMux I__656 (
            .O(N__4306),
            .I(N__4296));
    InMux I__655 (
            .O(N__4303),
            .I(N__4296));
    LocalMux I__654 (
            .O(N__4296),
            .I(\fsm_ctrl_inst1.counter_dinZ0Z_3 ));
    CascadeMux I__653 (
            .O(N__4293),
            .I(N__4289));
    InMux I__652 (
            .O(N__4292),
            .I(N__4275));
    InMux I__651 (
            .O(N__4289),
            .I(N__4275));
    InMux I__650 (
            .O(N__4288),
            .I(N__4275));
    InMux I__649 (
            .O(N__4287),
            .I(N__4275));
    InMux I__648 (
            .O(N__4286),
            .I(N__4275));
    LocalMux I__647 (
            .O(N__4275),
            .I(\fsm_ctrl_inst1.counter_dinZ0Z_1 ));
    InMux I__646 (
            .O(N__4272),
            .I(N__4264));
    InMux I__645 (
            .O(N__4271),
            .I(N__4255));
    InMux I__644 (
            .O(N__4270),
            .I(N__4255));
    InMux I__643 (
            .O(N__4269),
            .I(N__4255));
    InMux I__642 (
            .O(N__4268),
            .I(N__4255));
    InMux I__641 (
            .O(N__4267),
            .I(N__4252));
    LocalMux I__640 (
            .O(N__4264),
            .I(N__4247));
    LocalMux I__639 (
            .O(N__4255),
            .I(N__4247));
    LocalMux I__638 (
            .O(N__4252),
            .I(\fsm_ctrl_inst1.counter_dinZ0Z_0 ));
    Odrv4 I__637 (
            .O(N__4247),
            .I(\fsm_ctrl_inst1.counter_dinZ0Z_0 ));
    CascadeMux I__636 (
            .O(N__4242),
            .I(\fsm_ctrl_inst1.o2_cascade_ ));
    InMux I__635 (
            .O(N__4239),
            .I(N__4236));
    LocalMux I__634 (
            .O(N__4236),
            .I(\config_register_latched_dec_inst1.STATSRZ0Z_0 ));
    InMux I__633 (
            .O(N__4233),
            .I(N__4230));
    LocalMux I__632 (
            .O(N__4230),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_19 ));
    InMux I__631 (
            .O(N__4227),
            .I(N__4224));
    LocalMux I__630 (
            .O(N__4224),
            .I(N__4221));
    Odrv4 I__629 (
            .O(N__4221),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_20 ));
    CEMux I__628 (
            .O(N__4218),
            .I(N__4155));
    CEMux I__627 (
            .O(N__4217),
            .I(N__4155));
    CEMux I__626 (
            .O(N__4216),
            .I(N__4155));
    CEMux I__625 (
            .O(N__4215),
            .I(N__4155));
    CEMux I__624 (
            .O(N__4214),
            .I(N__4155));
    CEMux I__623 (
            .O(N__4213),
            .I(N__4155));
    CEMux I__622 (
            .O(N__4212),
            .I(N__4155));
    CEMux I__621 (
            .O(N__4211),
            .I(N__4155));
    CEMux I__620 (
            .O(N__4210),
            .I(N__4155));
    CEMux I__619 (
            .O(N__4209),
            .I(N__4155));
    CEMux I__618 (
            .O(N__4208),
            .I(N__4155));
    CEMux I__617 (
            .O(N__4207),
            .I(N__4155));
    CEMux I__616 (
            .O(N__4206),
            .I(N__4155));
    CEMux I__615 (
            .O(N__4205),
            .I(N__4155));
    CEMux I__614 (
            .O(N__4204),
            .I(N__4155));
    CEMux I__613 (
            .O(N__4203),
            .I(N__4155));
    CEMux I__612 (
            .O(N__4202),
            .I(N__4155));
    CEMux I__611 (
            .O(N__4201),
            .I(N__4155));
    CEMux I__610 (
            .O(N__4200),
            .I(N__4155));
    CEMux I__609 (
            .O(N__4199),
            .I(N__4155));
    CEMux I__608 (
            .O(N__4198),
            .I(N__4155));
    GlobalMux I__607 (
            .O(N__4155),
            .I(N__4152));
    gio2CtrlBuf I__606 (
            .O(N__4152),
            .I(\fsm_ctrl_inst1.current_state_i_g_0 ));
    IoInMux I__605 (
            .O(N__4149),
            .I(N__4146));
    LocalMux I__604 (
            .O(N__4146),
            .I(N__4143));
    IoSpan4Mux I__603 (
            .O(N__4143),
            .I(N__4140));
    Span4Mux_s3_h I__602 (
            .O(N__4140),
            .I(N__4137));
    Odrv4 I__601 (
            .O(N__4137),
            .I(SDO_signal_out_c));
    InMux I__600 (
            .O(N__4134),
            .I(N__4131));
    LocalMux I__599 (
            .O(N__4131),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_31 ));
    InMux I__598 (
            .O(N__4128),
            .I(N__4125));
    LocalMux I__597 (
            .O(N__4125),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_32 ));
    InMux I__596 (
            .O(N__4122),
            .I(N__4109));
    InMux I__595 (
            .O(N__4121),
            .I(N__4109));
    InMux I__594 (
            .O(N__4120),
            .I(N__4109));
    InMux I__593 (
            .O(N__4119),
            .I(N__4106));
    InMux I__592 (
            .O(N__4118),
            .I(N__4103));
    InMux I__591 (
            .O(N__4117),
            .I(N__4100));
    InMux I__590 (
            .O(N__4116),
            .I(N__4097));
    LocalMux I__589 (
            .O(N__4109),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_1 ));
    LocalMux I__588 (
            .O(N__4106),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_1 ));
    LocalMux I__587 (
            .O(N__4103),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_1 ));
    LocalMux I__586 (
            .O(N__4100),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_1 ));
    LocalMux I__585 (
            .O(N__4097),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_1 ));
    CascadeMux I__584 (
            .O(N__4086),
            .I(N__4081));
    CascadeMux I__583 (
            .O(N__4085),
            .I(N__4078));
    InMux I__582 (
            .O(N__4084),
            .I(N__4071));
    InMux I__581 (
            .O(N__4081),
            .I(N__4064));
    InMux I__580 (
            .O(N__4078),
            .I(N__4064));
    InMux I__579 (
            .O(N__4077),
            .I(N__4064));
    InMux I__578 (
            .O(N__4076),
            .I(N__4061));
    InMux I__577 (
            .O(N__4075),
            .I(N__4058));
    InMux I__576 (
            .O(N__4074),
            .I(N__4055));
    LocalMux I__575 (
            .O(N__4071),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_3 ));
    LocalMux I__574 (
            .O(N__4064),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_3 ));
    LocalMux I__573 (
            .O(N__4061),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_3 ));
    LocalMux I__572 (
            .O(N__4058),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_3 ));
    LocalMux I__571 (
            .O(N__4055),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_3 ));
    InMux I__570 (
            .O(N__4044),
            .I(N__4039));
    InMux I__569 (
            .O(N__4043),
            .I(N__4036));
    InMux I__568 (
            .O(N__4042),
            .I(N__4033));
    LocalMux I__567 (
            .O(N__4039),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_0 ));
    LocalMux I__566 (
            .O(N__4036),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_0 ));
    LocalMux I__565 (
            .O(N__4033),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_0 ));
    InMux I__564 (
            .O(N__4026),
            .I(N__4023));
    LocalMux I__563 (
            .O(N__4023),
            .I(\fsm_ctrl_inst1.current_state_RNO_2Z0Z_0 ));
    InMux I__562 (
            .O(N__4020),
            .I(N__4017));
    LocalMux I__561 (
            .O(N__4017),
            .I(\fsm_ctrl_inst1.g0_0_3_0 ));
    CascadeMux I__560 (
            .O(N__4014),
            .I(N__4007));
    CascadeMux I__559 (
            .O(N__4013),
            .I(N__4002));
    InMux I__558 (
            .O(N__4012),
            .I(N__3999));
    InMux I__557 (
            .O(N__4011),
            .I(N__3996));
    InMux I__556 (
            .O(N__4010),
            .I(N__3993));
    InMux I__555 (
            .O(N__4007),
            .I(N__3990));
    InMux I__554 (
            .O(N__4006),
            .I(N__3983));
    InMux I__553 (
            .O(N__4005),
            .I(N__3983));
    InMux I__552 (
            .O(N__4002),
            .I(N__3983));
    LocalMux I__551 (
            .O(N__3999),
            .I(\fsm_ctrl_inst1.counter_idleZ1Z_4 ));
    LocalMux I__550 (
            .O(N__3996),
            .I(\fsm_ctrl_inst1.counter_idleZ1Z_4 ));
    LocalMux I__549 (
            .O(N__3993),
            .I(\fsm_ctrl_inst1.counter_idleZ1Z_4 ));
    LocalMux I__548 (
            .O(N__3990),
            .I(\fsm_ctrl_inst1.counter_idleZ1Z_4 ));
    LocalMux I__547 (
            .O(N__3983),
            .I(\fsm_ctrl_inst1.counter_idleZ1Z_4 ));
    InMux I__546 (
            .O(N__3972),
            .I(N__3963));
    InMux I__545 (
            .O(N__3971),
            .I(N__3958));
    InMux I__544 (
            .O(N__3970),
            .I(N__3958));
    InMux I__543 (
            .O(N__3969),
            .I(N__3955));
    InMux I__542 (
            .O(N__3968),
            .I(N__3950));
    InMux I__541 (
            .O(N__3967),
            .I(N__3950));
    InMux I__540 (
            .O(N__3966),
            .I(N__3947));
    LocalMux I__539 (
            .O(N__3963),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_2 ));
    LocalMux I__538 (
            .O(N__3958),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_2 ));
    LocalMux I__537 (
            .O(N__3955),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_2 ));
    LocalMux I__536 (
            .O(N__3950),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_2 ));
    LocalMux I__535 (
            .O(N__3947),
            .I(\fsm_ctrl_inst1.counter_idleZ0Z_2 ));
    InMux I__534 (
            .O(N__3936),
            .I(N__3933));
    LocalMux I__533 (
            .O(N__3933),
            .I(\fsm_ctrl_inst1.g0_0_3 ));
    CascadeMux I__532 (
            .O(N__3930),
            .I(\fsm_ctrl_inst1.counter_din_RNO_0Z0Z_3_cascade_ ));
    CascadeMux I__531 (
            .O(N__3927),
            .I(\fsm_ctrl_inst1.current_state_RNO_3Z0Z_0_cascade_ ));
    InMux I__530 (
            .O(N__3924),
            .I(N__3921));
    LocalMux I__529 (
            .O(N__3921),
            .I(\fsm_ctrl_inst1.current_state_RNO_1Z0Z_0 ));
    InMux I__528 (
            .O(N__3918),
            .I(N__3915));
    LocalMux I__527 (
            .O(N__3915),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_23 ));
    InMux I__526 (
            .O(N__3912),
            .I(N__3909));
    LocalMux I__525 (
            .O(N__3909),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_24 ));
    InMux I__524 (
            .O(N__3906),
            .I(N__3903));
    LocalMux I__523 (
            .O(N__3903),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_45 ));
    InMux I__522 (
            .O(N__3900),
            .I(N__3897));
    LocalMux I__521 (
            .O(N__3897),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_46 ));
    InMux I__520 (
            .O(N__3894),
            .I(N__3891));
    LocalMux I__519 (
            .O(N__3891),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_27 ));
    InMux I__518 (
            .O(N__3888),
            .I(N__3885));
    LocalMux I__517 (
            .O(N__3885),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_28 ));
    InMux I__516 (
            .O(N__3882),
            .I(N__3879));
    LocalMux I__515 (
            .O(N__3879),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_33 ));
    InMux I__514 (
            .O(N__3876),
            .I(N__3873));
    LocalMux I__513 (
            .O(N__3873),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_29 ));
    InMux I__512 (
            .O(N__3870),
            .I(N__3867));
    LocalMux I__511 (
            .O(N__3867),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_34 ));
    InMux I__510 (
            .O(N__3864),
            .I(N__3861));
    LocalMux I__509 (
            .O(N__3861),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_30 ));
    InMux I__508 (
            .O(N__3858),
            .I(N__3855));
    LocalMux I__507 (
            .O(N__3855),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_35 ));
    InMux I__506 (
            .O(N__3852),
            .I(N__3849));
    LocalMux I__505 (
            .O(N__3849),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_36 ));
    InMux I__504 (
            .O(N__3846),
            .I(N__3843));
    LocalMux I__503 (
            .O(N__3843),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_26 ));
    InMux I__502 (
            .O(N__3840),
            .I(N__3837));
    LocalMux I__501 (
            .O(N__3837),
            .I(N__3834));
    Odrv4 I__500 (
            .O(N__3834),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_12 ));
    InMux I__499 (
            .O(N__3831),
            .I(N__3828));
    LocalMux I__498 (
            .O(N__3828),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_13 ));
    InMux I__497 (
            .O(N__3825),
            .I(N__3822));
    LocalMux I__496 (
            .O(N__3822),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_49 ));
    InMux I__495 (
            .O(N__3819),
            .I(N__3816));
    LocalMux I__494 (
            .O(N__3816),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_50 ));
    InMux I__493 (
            .O(N__3813),
            .I(N__3810));
    LocalMux I__492 (
            .O(N__3810),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_47 ));
    InMux I__491 (
            .O(N__3807),
            .I(N__3804));
    LocalMux I__490 (
            .O(N__3804),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_25 ));
    InMux I__489 (
            .O(N__3801),
            .I(N__3798));
    LocalMux I__488 (
            .O(N__3798),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_44 ));
    InMux I__487 (
            .O(N__3795),
            .I(N__3792));
    LocalMux I__486 (
            .O(N__3792),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_51 ));
    InMux I__485 (
            .O(N__3789),
            .I(N__3786));
    LocalMux I__484 (
            .O(N__3786),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_52 ));
    InMux I__483 (
            .O(N__3783),
            .I(N__3780));
    LocalMux I__482 (
            .O(N__3780),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_17 ));
    InMux I__481 (
            .O(N__3777),
            .I(N__3774));
    LocalMux I__480 (
            .O(N__3774),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_16 ));
    InMux I__479 (
            .O(N__3771),
            .I(N__3768));
    LocalMux I__478 (
            .O(N__3768),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_14 ));
    InMux I__477 (
            .O(N__3765),
            .I(N__3762));
    LocalMux I__476 (
            .O(N__3762),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_15 ));
    InMux I__475 (
            .O(N__3759),
            .I(N__3756));
    LocalMux I__474 (
            .O(N__3756),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_62 ));
    InMux I__473 (
            .O(N__3753),
            .I(N__3750));
    LocalMux I__472 (
            .O(N__3750),
            .I(N__3747));
    Odrv12 I__471 (
            .O(N__3747),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_63 ));
    InMux I__470 (
            .O(N__3744),
            .I(N__3741));
    LocalMux I__469 (
            .O(N__3741),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_21 ));
    InMux I__468 (
            .O(N__3738),
            .I(N__3735));
    LocalMux I__467 (
            .O(N__3735),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_22 ));
    InMux I__466 (
            .O(N__3732),
            .I(N__3729));
    LocalMux I__465 (
            .O(N__3729),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_48 ));
    InMux I__464 (
            .O(N__3726),
            .I(N__3723));
    LocalMux I__463 (
            .O(N__3723),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_65 ));
    InMux I__462 (
            .O(N__3720),
            .I(N__3717));
    LocalMux I__461 (
            .O(N__3717),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_66 ));
    InMux I__460 (
            .O(N__3714),
            .I(N__3711));
    LocalMux I__459 (
            .O(N__3711),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_68 ));
    InMux I__458 (
            .O(N__3708),
            .I(N__3705));
    LocalMux I__457 (
            .O(N__3705),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_69 ));
    InMux I__456 (
            .O(N__3702),
            .I(N__3699));
    LocalMux I__455 (
            .O(N__3699),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_70 ));
    InMux I__454 (
            .O(N__3696),
            .I(N__3693));
    LocalMux I__453 (
            .O(N__3693),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_73 ));
    InMux I__452 (
            .O(N__3690),
            .I(N__3687));
    LocalMux I__451 (
            .O(N__3687),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_74 ));
    InMux I__450 (
            .O(N__3684),
            .I(N__3681));
    LocalMux I__449 (
            .O(N__3681),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_71 ));
    InMux I__448 (
            .O(N__3678),
            .I(N__3675));
    LocalMux I__447 (
            .O(N__3675),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_72 ));
    InMux I__446 (
            .O(N__3672),
            .I(N__3669));
    LocalMux I__445 (
            .O(N__3669),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_18 ));
    CascadeMux I__444 (
            .O(N__3666),
            .I(\fsm_ctrl_inst1.counter_idle_RNO_1Z0Z_0_cascade_ ));
    CascadeMux I__443 (
            .O(N__3663),
            .I(\fsm_ctrl_inst1.counter_idlee_0_cascade_ ));
    InMux I__442 (
            .O(N__3660),
            .I(N__3657));
    LocalMux I__441 (
            .O(N__3657),
            .I(\fsm_ctrl_inst1.counter_idle_s_1 ));
    InMux I__440 (
            .O(N__3654),
            .I(N__3651));
    LocalMux I__439 (
            .O(N__3651),
            .I(\fsm_ctrl_inst1.g0_0_3_2 ));
    CascadeMux I__438 (
            .O(N__3648),
            .I(N__3645));
    InMux I__437 (
            .O(N__3645),
            .I(N__3642));
    LocalMux I__436 (
            .O(N__3642),
            .I(\fsm_ctrl_inst1.g0_0_2_2 ));
    InMux I__435 (
            .O(N__3639),
            .I(N__3631));
    InMux I__434 (
            .O(N__3638),
            .I(N__3631));
    InMux I__433 (
            .O(N__3637),
            .I(N__3626));
    InMux I__432 (
            .O(N__3636),
            .I(N__3626));
    LocalMux I__431 (
            .O(N__3631),
            .I(\fsm_ctrl_inst1.current_state_20_d_i ));
    LocalMux I__430 (
            .O(N__3626),
            .I(\fsm_ctrl_inst1.current_state_20_d_i ));
    InMux I__429 (
            .O(N__3621),
            .I(N__3618));
    LocalMux I__428 (
            .O(N__3618),
            .I(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_15 ));
    CascadeMux I__427 (
            .O(N__3615),
            .I(N__3612));
    InMux I__426 (
            .O(N__3612),
            .I(N__3609));
    LocalMux I__425 (
            .O(N__3609),
            .I(N__3606));
    Span4Mux_v I__424 (
            .O(N__3606),
            .I(N__3603));
    Odrv4 I__423 (
            .O(N__3603),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_87 ));
    InMux I__422 (
            .O(N__3600),
            .I(N__3597));
    LocalMux I__421 (
            .O(N__3597),
            .I(N__3594));
    Odrv4 I__420 (
            .O(N__3594),
            .I(CONSTANT_ONE_NET));
    InMux I__419 (
            .O(N__3591),
            .I(N__3588));
    LocalMux I__418 (
            .O(N__3588),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_67 ));
    InMux I__417 (
            .O(N__3585),
            .I(N__3582));
    LocalMux I__416 (
            .O(N__3582),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_64 ));
    CascadeMux I__415 (
            .O(N__3579),
            .I(\fsm_ctrl_inst1.g0_0_2_0_cascade_ ));
    InMux I__414 (
            .O(N__3576),
            .I(N__3573));
    LocalMux I__413 (
            .O(N__3573),
            .I(\fsm_ctrl_inst1.counter_idle_s_3 ));
    CascadeMux I__412 (
            .O(N__3570),
            .I(\fsm_ctrl_inst1.g0_0_2_cascade_ ));
    InMux I__411 (
            .O(N__3567),
            .I(N__3564));
    LocalMux I__410 (
            .O(N__3564),
            .I(\fsm_ctrl_inst1.counter_idle_s_4 ));
    InMux I__409 (
            .O(N__3561),
            .I(N__3558));
    LocalMux I__408 (
            .O(N__3558),
            .I(\fsm_ctrl_inst1.g0_0_3_1 ));
    InMux I__407 (
            .O(N__3555),
            .I(N__3552));
    LocalMux I__406 (
            .O(N__3552),
            .I(\fsm_ctrl_inst1.g0_0_2_1 ));
    CascadeMux I__405 (
            .O(N__3549),
            .I(\fsm_ctrl_inst1.current_state_20_d_i_cascade_ ));
    InMux I__404 (
            .O(N__3546),
            .I(N__3543));
    LocalMux I__403 (
            .O(N__3543),
            .I(\fsm_ctrl_inst1.counter_idle_s_2 ));
    CascadeMux I__402 (
            .O(N__3540),
            .I(\fsm_ctrl_inst1.N_93_0_cascade_ ));
    InMux I__401 (
            .O(N__3537),
            .I(N__3534));
    LocalMux I__400 (
            .O(N__3534),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_3 ));
    InMux I__399 (
            .O(N__3531),
            .I(N__3528));
    LocalMux I__398 (
            .O(N__3528),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_1 ));
    InMux I__397 (
            .O(N__3525),
            .I(N__3522));
    LocalMux I__396 (
            .O(N__3522),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_2 ));
    InMux I__395 (
            .O(N__3519),
            .I(N__3516));
    LocalMux I__394 (
            .O(N__3516),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_38 ));
    InMux I__393 (
            .O(N__3513),
            .I(N__3510));
    LocalMux I__392 (
            .O(N__3510),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_39 ));
    InMux I__391 (
            .O(N__3507),
            .I(N__3504));
    LocalMux I__390 (
            .O(N__3504),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_0 ));
    InMux I__389 (
            .O(N__3501),
            .I(N__3498));
    LocalMux I__388 (
            .O(N__3498),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_40 ));
    InMux I__387 (
            .O(N__3495),
            .I(N__3492));
    LocalMux I__386 (
            .O(N__3492),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_41 ));
    InMux I__385 (
            .O(N__3489),
            .I(N__3486));
    LocalMux I__384 (
            .O(N__3486),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_43 ));
    InMux I__383 (
            .O(N__3483),
            .I(N__3480));
    LocalMux I__382 (
            .O(N__3480),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_80 ));
    InMux I__381 (
            .O(N__3477),
            .I(N__3474));
    LocalMux I__380 (
            .O(N__3474),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_4 ));
    InMux I__379 (
            .O(N__3471),
            .I(N__3468));
    LocalMux I__378 (
            .O(N__3468),
            .I(N__3465));
    Odrv12 I__377 (
            .O(N__3465),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_5 ));
    InMux I__376 (
            .O(N__3462),
            .I(N__3459));
    LocalMux I__375 (
            .O(N__3459),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_53 ));
    InMux I__374 (
            .O(N__3456),
            .I(N__3453));
    LocalMux I__373 (
            .O(N__3453),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_37 ));
    InMux I__372 (
            .O(N__3450),
            .I(N__3447));
    LocalMux I__371 (
            .O(N__3447),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_81 ));
    InMux I__370 (
            .O(N__3444),
            .I(N__3441));
    LocalMux I__369 (
            .O(N__3441),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_82 ));
    InMux I__368 (
            .O(N__3438),
            .I(N__3435));
    LocalMux I__367 (
            .O(N__3435),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_75 ));
    InMux I__366 (
            .O(N__3432),
            .I(N__3429));
    LocalMux I__365 (
            .O(N__3429),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_76 ));
    InMux I__364 (
            .O(N__3426),
            .I(N__3423));
    LocalMux I__363 (
            .O(N__3423),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_77 ));
    InMux I__362 (
            .O(N__3420),
            .I(N__3417));
    LocalMux I__361 (
            .O(N__3417),
            .I(N__3414));
    Odrv4 I__360 (
            .O(N__3414),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_11 ));
    InMux I__359 (
            .O(N__3411),
            .I(N__3408));
    LocalMux I__358 (
            .O(N__3408),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_54 ));
    InMux I__357 (
            .O(N__3405),
            .I(N__3402));
    LocalMux I__356 (
            .O(N__3402),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_60 ));
    InMux I__355 (
            .O(N__3399),
            .I(N__3396));
    LocalMux I__354 (
            .O(N__3396),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_61 ));
    InMux I__353 (
            .O(N__3393),
            .I(N__3390));
    LocalMux I__352 (
            .O(N__3390),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_78 ));
    InMux I__351 (
            .O(N__3387),
            .I(N__3384));
    LocalMux I__350 (
            .O(N__3384),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_79 ));
    InMux I__349 (
            .O(N__3381),
            .I(N__3378));
    LocalMux I__348 (
            .O(N__3378),
            .I(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_9 ));
    InMux I__347 (
            .O(N__3375),
            .I(N__3372));
    LocalMux I__346 (
            .O(N__3372),
            .I(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_6 ));
    InMux I__345 (
            .O(N__3369),
            .I(N__3366));
    LocalMux I__344 (
            .O(N__3366),
            .I(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_7 ));
    InMux I__343 (
            .O(N__3363),
            .I(N__3360));
    LocalMux I__342 (
            .O(N__3360),
            .I(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_8 ));
    InMux I__341 (
            .O(N__3357),
            .I(N__3354));
    LocalMux I__340 (
            .O(N__3354),
            .I(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_12 ));
    InMux I__339 (
            .O(N__3351),
            .I(N__3348));
    LocalMux I__338 (
            .O(N__3348),
            .I(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_10 ));
    InMux I__337 (
            .O(N__3345),
            .I(N__3342));
    LocalMux I__336 (
            .O(N__3342),
            .I(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_11 ));
    InMux I__335 (
            .O(N__3339),
            .I(N__3336));
    LocalMux I__334 (
            .O(N__3336),
            .I(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_13 ));
    InMux I__333 (
            .O(N__3333),
            .I(N__3330));
    LocalMux I__332 (
            .O(N__3330),
            .I(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_14 ));
    CEMux I__331 (
            .O(N__3327),
            .I(N__3322));
    CEMux I__330 (
            .O(N__3326),
            .I(N__3319));
    CEMux I__329 (
            .O(N__3325),
            .I(N__3316));
    LocalMux I__328 (
            .O(N__3322),
            .I(N__3313));
    LocalMux I__327 (
            .O(N__3319),
            .I(N__3308));
    LocalMux I__326 (
            .O(N__3316),
            .I(N__3308));
    Odrv4 I__325 (
            .O(N__3313),
            .I(\fsm_ctrl_inst1.current_state_i_1 ));
    Odrv4 I__324 (
            .O(N__3308),
            .I(\fsm_ctrl_inst1.current_state_i_1 ));
    InMux I__323 (
            .O(N__3303),
            .I(N__3300));
    LocalMux I__322 (
            .O(N__3300),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_42 ));
    InMux I__321 (
            .O(N__3297),
            .I(\fsm_ctrl_inst1.counter_idle_cry_0 ));
    InMux I__320 (
            .O(N__3294),
            .I(\fsm_ctrl_inst1.counter_idle_cry_1 ));
    InMux I__319 (
            .O(N__3291),
            .I(\fsm_ctrl_inst1.counter_idle_cry_2 ));
    InMux I__318 (
            .O(N__3288),
            .I(\fsm_ctrl_inst1.counter_idle_cry_3 ));
    InMux I__317 (
            .O(N__3285),
            .I(N__3282));
    LocalMux I__316 (
            .O(N__3282),
            .I(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_3 ));
    InMux I__315 (
            .O(N__3279),
            .I(N__3276));
    LocalMux I__314 (
            .O(N__3276),
            .I(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_4 ));
    InMux I__313 (
            .O(N__3273),
            .I(N__3270));
    LocalMux I__312 (
            .O(N__3270),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_56 ));
    InMux I__311 (
            .O(N__3267),
            .I(N__3264));
    LocalMux I__310 (
            .O(N__3264),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_59 ));
    InMux I__309 (
            .O(N__3261),
            .I(N__3258));
    LocalMux I__308 (
            .O(N__3258),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_55 ));
    InMux I__307 (
            .O(N__3255),
            .I(N__3252));
    LocalMux I__306 (
            .O(N__3252),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_7 ));
    InMux I__305 (
            .O(N__3249),
            .I(N__3246));
    LocalMux I__304 (
            .O(N__3246),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_8 ));
    InMux I__303 (
            .O(N__3243),
            .I(N__3240));
    LocalMux I__302 (
            .O(N__3240),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_9 ));
    InMux I__301 (
            .O(N__3237),
            .I(N__3234));
    LocalMux I__300 (
            .O(N__3234),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_10 ));
    InMux I__299 (
            .O(N__3231),
            .I(N__3228));
    LocalMux I__298 (
            .O(N__3228),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_83 ));
    InMux I__297 (
            .O(N__3225),
            .I(N__3222));
    LocalMux I__296 (
            .O(N__3222),
            .I(N__3219));
    Odrv4 I__295 (
            .O(N__3219),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_84 ));
    InMux I__294 (
            .O(N__3216),
            .I(N__3213));
    LocalMux I__293 (
            .O(N__3213),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_85 ));
    InMux I__292 (
            .O(N__3210),
            .I(N__3207));
    LocalMux I__291 (
            .O(N__3207),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_86 ));
    InMux I__290 (
            .O(N__3204),
            .I(N__3201));
    LocalMux I__289 (
            .O(N__3201),
            .I(N__3198));
    Odrv4 I__288 (
            .O(N__3198),
            .I(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_1 ));
    InMux I__287 (
            .O(N__3195),
            .I(N__3192));
    LocalMux I__286 (
            .O(N__3192),
            .I(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_2 ));
    InMux I__285 (
            .O(N__3189),
            .I(N__3186));
    LocalMux I__284 (
            .O(N__3186),
            .I(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_5 ));
    InMux I__283 (
            .O(N__3183),
            .I(N__3180));
    LocalMux I__282 (
            .O(N__3180),
            .I(N__3177));
    Span4Mux_v I__281 (
            .O(N__3177),
            .I(N__3174));
    Odrv4 I__280 (
            .O(N__3174),
            .I(RST_N_c));
    IoInMux I__279 (
            .O(N__3171),
            .I(N__3168));
    LocalMux I__278 (
            .O(N__3168),
            .I(N__3165));
    Span12Mux_s0_h I__277 (
            .O(N__3165),
            .I(N__3162));
    Odrv12 I__276 (
            .O(N__3162),
            .I(RST_N_c_i));
    IoInMux I__275 (
            .O(N__3159),
            .I(N__3156));
    LocalMux I__274 (
            .O(N__3156),
            .I(\fsm_ctrl_inst1.current_state_i_0 ));
    InMux I__273 (
            .O(N__3153),
            .I(N__3150));
    LocalMux I__272 (
            .O(N__3150),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_58 ));
    InMux I__271 (
            .O(N__3147),
            .I(N__3144));
    LocalMux I__270 (
            .O(N__3144),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_57 ));
    InMux I__269 (
            .O(N__3141),
            .I(N__3138));
    LocalMux I__268 (
            .O(N__3138),
            .I(\fsm_ctrl_inst1.bit_sequence_statZ0Z_6 ));
    InMux I__267 (
            .O(N__3135),
            .I(N__3132));
    LocalMux I__266 (
            .O(N__3132),
            .I(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_0 ));
    defparam IN_MUX_bfv_3_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_20_0_));
    ICE_GB N_218_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4608),
            .GLOBALBUFFEROUTPUT(N_218_g));
    ICE_GB \fsm_ctrl_inst1.current_state_RNI1GR8_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__3159),
            .GLOBALBUFFEROUTPUT(\fsm_ctrl_inst1.current_state_i_g_0 ));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB RST_N_ibuf_RNIBJGC_0 (
            .USERSIGNALTOGLOBALBUFFER(N__3171),
            .GLOBALBUFFEROUTPUT(RST_N_c_i_g));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam RST_N_ibuf_RNIBJGC_LC_1_6_2.C_ON=1'b0;
    defparam RST_N_ibuf_RNIBJGC_LC_1_6_2.SEQ_MODE=4'b0000;
    defparam RST_N_ibuf_RNIBJGC_LC_1_6_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 RST_N_ibuf_RNIBJGC_LC_1_6_2 (
            .in0(N__3183),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RST_N_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.current_state_RNI1GR8_0_LC_1_17_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.current_state_RNI1GR8_0_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.current_state_RNI1GR8_0_LC_1_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \fsm_ctrl_inst1.current_state_RNI1GR8_0_LC_1_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4596),
            .lcout(\fsm_ctrl_inst1.current_state_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_58_LC_2_16_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_58_LC_2_16_0 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_58_LC_2_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_58_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__3147),
            .in2(_gnd_net_),
            .in3(N__5036),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6121),
            .ce(N__4200),
            .sr(N__5801));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_59_LC_2_17_2 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_59_LC_2_17_2 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_59_LC_2_17_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_59_LC_2_17_2  (
            .in0(N__5055),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3153),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6119),
            .ce(N__4198),
            .sr(N__5802));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_57_LC_2_17_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_57_LC_2_17_3 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_57_LC_2_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_57_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(N__3273),
            .in2(_gnd_net_),
            .in3(N__5054),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6119),
            .ce(N__4198),
            .sr(N__5802));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_7_LC_2_18_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_7_LC_2_18_5 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_7_LC_2_18_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_7_LC_2_18_5  (
            .in0(_gnd_net_),
            .in1(N__3141),
            .in2(_gnd_net_),
            .in3(N__4984),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6122),
            .ce(N__4201),
            .sr(N__5804));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_6_LC_2_18_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_6_LC_2_18_7 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_6_LC_2_18_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_6_LC_2_18_7  (
            .in0(_gnd_net_),
            .in1(N__3471),
            .in2(_gnd_net_),
            .in3(N__4983),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6122),
            .ce(N__4201),
            .sr(N__5804));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_84_LC_2_19_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_84_LC_2_19_4 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_84_LC_2_19_4 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_84_LC_2_19_4  (
            .in0(_gnd_net_),
            .in1(N__3231),
            .in2(_gnd_net_),
            .in3(N__4972),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6124),
            .ce(N__4203),
            .sr(N__5807));
    defparam \fsm_ctrl_inst1.bit_sequence_din_1_LC_2_20_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_din_1_LC_2_20_3 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_din_1_LC_2_20_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_din_1_LC_2_20_3  (
            .in0(N__4588),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3135),
            .lcout(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6127),
            .ce(N__3325),
            .sr(N__5811));
    defparam \fsm_ctrl_inst1.bit_sequence_din_0_LC_2_20_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_din_0_LC_2_20_4 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_din_0_LC_2_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_din_0_LC_2_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4589),
            .lcout(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6127),
            .ce(N__3325),
            .sr(N__5811));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_85_LC_2_21_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_85_LC_2_21_3 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_85_LC_2_21_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_85_LC_2_21_3  (
            .in0(_gnd_net_),
            .in1(N__3225),
            .in2(_gnd_net_),
            .in3(N__4962),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6131),
            .ce(N__4209),
            .sr(N__5816));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_86_LC_2_21_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_86_LC_2_21_4 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_86_LC_2_21_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_86_LC_2_21_4  (
            .in0(N__4963),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3216),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6131),
            .ce(N__4209),
            .sr(N__5816));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_87_LC_2_21_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_87_LC_2_21_5 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_87_LC_2_21_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_87_LC_2_21_5  (
            .in0(_gnd_net_),
            .in1(N__3210),
            .in2(_gnd_net_),
            .in3(N__4964),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6131),
            .ce(N__4209),
            .sr(N__5816));
    defparam \fsm_ctrl_inst1.current_state_RNI2HR8_1_LC_2_21_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.current_state_RNI2HR8_1_LC_2_21_7 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.current_state_RNI2HR8_1_LC_2_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \fsm_ctrl_inst1.current_state_RNI2HR8_1_LC_2_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4961),
            .lcout(\fsm_ctrl_inst1.current_state_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.bit_sequence_din_3_LC_2_22_1 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_din_3_LC_2_22_1 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_din_3_LC_2_22_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_din_3_LC_2_22_1  (
            .in0(_gnd_net_),
            .in1(N__3195),
            .in2(_gnd_net_),
            .in3(N__4591),
            .lcout(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6136),
            .ce(N__3326),
            .sr(N__5820));
    defparam \fsm_ctrl_inst1.bit_sequence_din_5_LC_2_22_2 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_din_5_LC_2_22_2 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_din_5_LC_2_22_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_din_5_LC_2_22_2  (
            .in0(N__4595),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3279),
            .lcout(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6136),
            .ce(N__3326),
            .sr(N__5820));
    defparam \fsm_ctrl_inst1.bit_sequence_din_10_LC_2_22_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_din_10_LC_2_22_3 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_din_10_LC_2_22_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_din_10_LC_2_22_3  (
            .in0(_gnd_net_),
            .in1(N__3381),
            .in2(_gnd_net_),
            .in3(N__4590),
            .lcout(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6136),
            .ce(N__3326),
            .sr(N__5820));
    defparam \fsm_ctrl_inst1.bit_sequence_din_2_LC_2_22_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_din_2_LC_2_22_4 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_din_2_LC_2_22_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_din_2_LC_2_22_4  (
            .in0(N__4594),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3204),
            .lcout(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6136),
            .ce(N__3326),
            .sr(N__5820));
    defparam \fsm_ctrl_inst1.bit_sequence_din_6_LC_2_22_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_din_6_LC_2_22_5 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_din_6_LC_2_22_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_din_6_LC_2_22_5  (
            .in0(_gnd_net_),
            .in1(N__3189),
            .in2(_gnd_net_),
            .in3(N__4593),
            .lcout(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6136),
            .ce(N__3326),
            .sr(N__5820));
    defparam \fsm_ctrl_inst1.bit_sequence_din_4_LC_2_22_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_din_4_LC_2_22_7 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_din_4_LC_2_22_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_din_4_LC_2_22_7  (
            .in0(_gnd_net_),
            .in1(N__3285),
            .in2(_gnd_net_),
            .in3(N__4592),
            .lcout(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6136),
            .ce(N__3326),
            .sr(N__5820));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_56_LC_3_17_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_56_LC_3_17_5 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_56_LC_3_17_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_56_LC_3_17_5  (
            .in0(_gnd_net_),
            .in1(N__3261),
            .in2(_gnd_net_),
            .in3(N__5038),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6120),
            .ce(N__4199),
            .sr(N__5805));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_60_LC_3_17_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_60_LC_3_17_6 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_60_LC_3_17_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_60_LC_3_17_6  (
            .in0(N__5039),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3267),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6120),
            .ce(N__4199),
            .sr(N__5805));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_55_LC_3_17_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_55_LC_3_17_7 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_55_LC_3_17_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_55_LC_3_17_7  (
            .in0(_gnd_net_),
            .in1(N__3411),
            .in2(_gnd_net_),
            .in3(N__5037),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6120),
            .ce(N__4199),
            .sr(N__5805));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_8_LC_3_18_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_8_LC_3_18_0 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_8_LC_3_18_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_8_LC_3_18_0  (
            .in0(N__4970),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3255),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6125),
            .ce(N__4204),
            .sr(N__5808));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_10_LC_3_18_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_10_LC_3_18_3 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_10_LC_3_18_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_10_LC_3_18_3  (
            .in0(_gnd_net_),
            .in1(N__3243),
            .in2(_gnd_net_),
            .in3(N__4967),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6125),
            .ce(N__4204),
            .sr(N__5808));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_9_LC_3_18_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_9_LC_3_18_5 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_9_LC_3_18_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_9_LC_3_18_5  (
            .in0(_gnd_net_),
            .in1(N__3249),
            .in2(_gnd_net_),
            .in3(N__4971),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6125),
            .ce(N__4204),
            .sr(N__5808));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_11_LC_3_18_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_11_LC_3_18_6 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_11_LC_3_18_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_11_LC_3_18_6  (
            .in0(N__4968),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3237),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6125),
            .ce(N__4204),
            .sr(N__5808));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_83_LC_3_18_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_83_LC_3_18_7 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_83_LC_3_18_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_83_LC_3_18_7  (
            .in0(_gnd_net_),
            .in1(N__3444),
            .in2(_gnd_net_),
            .in3(N__4969),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6125),
            .ce(N__4204),
            .sr(N__5808));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_42_LC_3_19_2 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_42_LC_3_19_2 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_42_LC_3_19_2 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_42_LC_3_19_2  (
            .in0(N__3495),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4965),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6128),
            .ce(N__4206),
            .sr(N__5812));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_43_LC_3_19_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_43_LC_3_19_4 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_43_LC_3_19_4 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_43_LC_3_19_4  (
            .in0(_gnd_net_),
            .in1(N__3303),
            .in2(_gnd_net_),
            .in3(N__4966),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6128),
            .ce(N__4206),
            .sr(N__5812));
    defparam \fsm_ctrl_inst1.counter_idle_cry_c_0_LC_3_20_0 .C_ON=1'b1;
    defparam \fsm_ctrl_inst1.counter_idle_cry_c_0_LC_3_20_0 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.counter_idle_cry_c_0_LC_3_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_cry_c_0_LC_3_20_0  (
            .in0(_gnd_net_),
            .in1(N__4042),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_20_0_),
            .carryout(\fsm_ctrl_inst1.counter_idle_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_idle_RNO_0_1_LC_3_20_1 .C_ON=1'b1;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_0_1_LC_3_20_1 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_0_1_LC_3_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_RNO_0_1_LC_3_20_1  (
            .in0(_gnd_net_),
            .in1(N__4116),
            .in2(_gnd_net_),
            .in3(N__3297),
            .lcout(\fsm_ctrl_inst1.counter_idle_s_1 ),
            .ltout(),
            .carryin(\fsm_ctrl_inst1.counter_idle_cry_0 ),
            .carryout(\fsm_ctrl_inst1.counter_idle_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_idle_RNO_0_2_LC_3_20_2 .C_ON=1'b1;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_0_2_LC_3_20_2 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_0_2_LC_3_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_RNO_0_2_LC_3_20_2  (
            .in0(_gnd_net_),
            .in1(N__3966),
            .in2(_gnd_net_),
            .in3(N__3294),
            .lcout(\fsm_ctrl_inst1.counter_idle_s_2 ),
            .ltout(),
            .carryin(\fsm_ctrl_inst1.counter_idle_cry_1 ),
            .carryout(\fsm_ctrl_inst1.counter_idle_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_idle_RNO_0_3_LC_3_20_3 .C_ON=1'b1;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_0_3_LC_3_20_3 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_0_3_LC_3_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_RNO_0_3_LC_3_20_3  (
            .in0(_gnd_net_),
            .in1(N__4075),
            .in2(_gnd_net_),
            .in3(N__3291),
            .lcout(\fsm_ctrl_inst1.counter_idle_s_3 ),
            .ltout(),
            .carryin(\fsm_ctrl_inst1.counter_idle_cry_2 ),
            .carryout(\fsm_ctrl_inst1.counter_idle_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_idle_RNO_0_4_LC_3_20_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_0_4_LC_3_20_4 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_0_4_LC_3_20_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_RNO_0_4_LC_3_20_4  (
            .in0(_gnd_net_),
            .in1(N__4010),
            .in2(_gnd_net_),
            .in3(N__3288),
            .lcout(\fsm_ctrl_inst1.counter_idle_s_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_idle_RNO_2_1_LC_3_21_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_2_1_LC_3_21_0 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_2_1_LC_3_21_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_RNO_2_1_LC_3_21_0  (
            .in0(N__4012),
            .in1(N__3972),
            .in2(N__4960),
            .in3(N__4543),
            .lcout(\fsm_ctrl_inst1.g0_0_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_din_0_LC_3_21_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_din_0_LC_3_21_4 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.counter_din_0_LC_3_21_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fsm_ctrl_inst1.counter_din_0_LC_3_21_4  (
            .in0(_gnd_net_),
            .in1(N__4267),
            .in2(_gnd_net_),
            .in3(N__4544),
            .lcout(\fsm_ctrl_inst1.counter_dinZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6137),
            .ce(),
            .sr(N__5821));
    defparam \fsm_ctrl_inst1.counter_idle_RNO_1_1_LC_3_21_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_1_1_LC_3_21_6 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_1_1_LC_3_21_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_RNO_1_1_LC_3_21_6  (
            .in0(_gnd_net_),
            .in1(N__4084),
            .in2(_gnd_net_),
            .in3(N__4119),
            .lcout(\fsm_ctrl_inst1.g0_0_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.bit_sequence_din_9_LC_3_22_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_din_9_LC_3_22_0 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_din_9_LC_3_22_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_din_9_LC_3_22_0  (
            .in0(_gnd_net_),
            .in1(N__4548),
            .in2(_gnd_net_),
            .in3(N__3363),
            .lcout(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6141),
            .ce(N__3327),
            .sr(N__5826));
    defparam \fsm_ctrl_inst1.bit_sequence_din_12_LC_3_22_1 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_din_12_LC_3_22_1 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_din_12_LC_3_22_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_din_12_LC_3_22_1  (
            .in0(N__4549),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3345),
            .lcout(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6141),
            .ce(N__3327),
            .sr(N__5826));
    defparam \fsm_ctrl_inst1.bit_sequence_din_7_LC_3_22_2 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_din_7_LC_3_22_2 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_din_7_LC_3_22_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_din_7_LC_3_22_2  (
            .in0(_gnd_net_),
            .in1(N__4547),
            .in2(_gnd_net_),
            .in3(N__3375),
            .lcout(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6141),
            .ce(N__3327),
            .sr(N__5826));
    defparam \fsm_ctrl_inst1.bit_sequence_din_8_LC_3_22_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_din_8_LC_3_22_3 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_din_8_LC_3_22_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_din_8_LC_3_22_3  (
            .in0(N__4552),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3369),
            .lcout(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6141),
            .ce(N__3327),
            .sr(N__5826));
    defparam \fsm_ctrl_inst1.bit_sequence_din_13_LC_3_22_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_din_13_LC_3_22_4 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_din_13_LC_3_22_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_din_13_LC_3_22_4  (
            .in0(_gnd_net_),
            .in1(N__4546),
            .in2(_gnd_net_),
            .in3(N__3357),
            .lcout(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6141),
            .ce(N__3327),
            .sr(N__5826));
    defparam \fsm_ctrl_inst1.bit_sequence_din_15_LC_3_22_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_din_15_LC_3_22_5 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_din_15_LC_3_22_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_din_15_LC_3_22_5  (
            .in0(N__4551),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3333),
            .lcout(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6141),
            .ce(N__3327),
            .sr(N__5826));
    defparam \fsm_ctrl_inst1.bit_sequence_din_11_LC_3_22_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_din_11_LC_3_22_6 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_din_11_LC_3_22_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_din_11_LC_3_22_6  (
            .in0(_gnd_net_),
            .in1(N__4545),
            .in2(_gnd_net_),
            .in3(N__3351),
            .lcout(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6141),
            .ce(N__3327),
            .sr(N__5826));
    defparam \fsm_ctrl_inst1.bit_sequence_din_14_LC_3_22_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_din_14_LC_3_22_7 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_din_14_LC_3_22_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_din_14_LC_3_22_7  (
            .in0(N__4550),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3339),
            .lcout(\fsm_ctrl_inst1.bit_sequence_dinZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6141),
            .ce(N__3327),
            .sr(N__5826));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_75_LC_4_15_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_75_LC_4_15_0 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_75_LC_4_15_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_75_LC_4_15_0  (
            .in0(N__5022),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3690),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6132),
            .ce(N__4210),
            .sr(N__5809));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_76_LC_4_15_1 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_76_LC_4_15_1 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_76_LC_4_15_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_76_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(N__3438),
            .in2(_gnd_net_),
            .in3(N__5023),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6132),
            .ce(N__4210),
            .sr(N__5809));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_77_LC_4_15_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_77_LC_4_15_4 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_77_LC_4_15_4 .LUT_INIT=16'b1101110111011101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_77_LC_4_15_4  (
            .in0(N__5024),
            .in1(N__3432),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6132),
            .ce(N__4210),
            .sr(N__5809));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_78_LC_4_16_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_78_LC_4_16_3 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_78_LC_4_16_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_78_LC_4_16_3  (
            .in0(N__5011),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3426),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6129),
            .ce(N__4207),
            .sr(N__5803));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_12_LC_4_16_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_12_LC_4_16_6 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_12_LC_4_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_12_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(N__3420),
            .in2(_gnd_net_),
            .in3(N__5010),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6129),
            .ce(N__4207),
            .sr(N__5803));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_54_LC_4_17_1 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_54_LC_4_17_1 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_54_LC_4_17_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_54_LC_4_17_1  (
            .in0(_gnd_net_),
            .in1(N__3462),
            .in2(_gnd_net_),
            .in3(N__5000),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6123),
            .ce(N__4202),
            .sr(N__5810));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_62_LC_4_17_2 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_62_LC_4_17_2 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_62_LC_4_17_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_62_LC_4_17_2  (
            .in0(N__5002),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3399),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6123),
            .ce(N__4202),
            .sr(N__5810));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_80_LC_4_17_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_80_LC_4_17_4 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_80_LC_4_17_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_80_LC_4_17_4  (
            .in0(N__5004),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3387),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6123),
            .ce(N__4202),
            .sr(N__5810));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_61_LC_4_17_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_61_LC_4_17_5 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_61_LC_4_17_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_61_LC_4_17_5  (
            .in0(_gnd_net_),
            .in1(N__3405),
            .in2(_gnd_net_),
            .in3(N__5001),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6123),
            .ce(N__4202),
            .sr(N__5810));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_79_LC_4_17_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_79_LC_4_17_6 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_79_LC_4_17_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_79_LC_4_17_6  (
            .in0(N__5003),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3393),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6123),
            .ce(N__4202),
            .sr(N__5810));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_4_LC_4_18_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_4_LC_4_18_0 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_4_LC_4_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_4_LC_4_18_0  (
            .in0(_gnd_net_),
            .in1(N__3537),
            .in2(_gnd_net_),
            .in3(N__4988),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6130),
            .ce(N__4208),
            .sr(N__5813));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_81_LC_4_18_1 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_81_LC_4_18_1 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_81_LC_4_18_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_81_LC_4_18_1  (
            .in0(N__4991),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3483),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6130),
            .ce(N__4208),
            .sr(N__5813));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_37_LC_4_18_2 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_37_LC_4_18_2 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_37_LC_4_18_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_37_LC_4_18_2  (
            .in0(N__3852),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4985),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6130),
            .ce(N__4208),
            .sr(N__5813));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_5_LC_4_18_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_5_LC_4_18_3 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_5_LC_4_18_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_5_LC_4_18_3  (
            .in0(N__4990),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3477),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6130),
            .ce(N__4208),
            .sr(N__5813));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_48_LC_4_18_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_48_LC_4_18_4 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_48_LC_4_18_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_48_LC_4_18_4  (
            .in0(_gnd_net_),
            .in1(N__3813),
            .in2(_gnd_net_),
            .in3(N__4987),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6130),
            .ce(N__4208),
            .sr(N__5813));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_53_LC_4_18_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_53_LC_4_18_5 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_53_LC_4_18_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_53_LC_4_18_5  (
            .in0(N__4989),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3789),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6130),
            .ce(N__4208),
            .sr(N__5813));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_38_LC_4_18_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_38_LC_4_18_6 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_38_LC_4_18_6 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_38_LC_4_18_6  (
            .in0(_gnd_net_),
            .in1(N__3456),
            .in2(_gnd_net_),
            .in3(N__4986),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6130),
            .ce(N__4208),
            .sr(N__5813));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_82_LC_4_18_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_82_LC_4_18_7 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_82_LC_4_18_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_82_LC_4_18_7  (
            .in0(N__4992),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3450),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6130),
            .ce(N__4208),
            .sr(N__5813));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_40_LC_4_19_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_40_LC_4_19_0 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_40_LC_4_19_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_40_LC_4_19_0  (
            .in0(N__4858),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3513),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6133),
            .ce(N__4211),
            .sr(N__5817));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_1_LC_4_19_1 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_1_LC_4_19_1 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_1_LC_4_19_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_1_LC_4_19_1  (
            .in0(_gnd_net_),
            .in1(N__3507),
            .in2(_gnd_net_),
            .in3(N__4854),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6133),
            .ce(N__4211),
            .sr(N__5817));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_3_LC_4_19_2 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_3_LC_4_19_2 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_3_LC_4_19_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_3_LC_4_19_2  (
            .in0(N__4857),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3525),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6133),
            .ce(N__4211),
            .sr(N__5817));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_2_LC_4_19_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_2_LC_4_19_3 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_2_LC_4_19_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_2_LC_4_19_3  (
            .in0(_gnd_net_),
            .in1(N__3531),
            .in2(_gnd_net_),
            .in3(N__4855),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6133),
            .ce(N__4211),
            .sr(N__5817));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_39_LC_4_19_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_39_LC_4_19_4 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_39_LC_4_19_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_39_LC_4_19_4  (
            .in0(N__4856),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3519),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6133),
            .ce(N__4211),
            .sr(N__5817));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_0_LC_4_19_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_0_LC_4_19_5 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_0_LC_4_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_0_LC_4_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4853),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6133),
            .ce(N__4211),
            .sr(N__5817));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_41_LC_4_19_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_41_LC_4_19_6 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_41_LC_4_19_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_41_LC_4_19_6  (
            .in0(N__4859),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3501),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6133),
            .ce(N__4211),
            .sr(N__5817));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_44_LC_4_19_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_44_LC_4_19_7 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_44_LC_4_19_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_44_LC_4_19_7  (
            .in0(_gnd_net_),
            .in1(N__3489),
            .in2(_gnd_net_),
            .in3(N__4860),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6133),
            .ce(N__4211),
            .sr(N__5817));
    defparam \fsm_ctrl_inst1.counter_idle_RNO_2_2_LC_4_20_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_2_2_LC_4_20_0 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_2_2_LC_4_20_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_RNO_2_2_LC_4_20_0  (
            .in0(N__4011),
            .in1(N__4542),
            .in2(N__4808),
            .in3(N__3969),
            .lcout(\fsm_ctrl_inst1.g0_0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_idle_RNO_1_2_LC_4_20_1 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_1_2_LC_4_20_1 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_1_2_LC_4_20_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_RNO_1_2_LC_4_20_1  (
            .in0(_gnd_net_),
            .in1(N__4077),
            .in2(_gnd_net_),
            .in3(N__4120),
            .lcout(\fsm_ctrl_inst1.g0_0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_idle_RNO_1_3_LC_4_20_2 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_1_3_LC_4_20_2 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_1_3_LC_4_20_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_RNO_1_3_LC_4_20_2  (
            .in0(N__4121),
            .in1(_gnd_net_),
            .in2(N__4085),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\fsm_ctrl_inst1.g0_0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_idle_3_LC_4_20_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_idle_3_LC_4_20_3 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.counter_idle_3_LC_4_20_3 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_3_LC_4_20_3  (
            .in0(N__4020),
            .in1(N__3636),
            .in2(N__3579),
            .in3(N__3576),
            .lcout(\fsm_ctrl_inst1.counter_idleZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6138),
            .ce(),
            .sr(N__5822));
    defparam \fsm_ctrl_inst1.counter_idle_RNO_1_4_LC_4_20_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_1_4_LC_4_20_4 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_1_4_LC_4_20_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_RNO_1_4_LC_4_20_4  (
            .in0(N__4122),
            .in1(_gnd_net_),
            .in2(N__4086),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\fsm_ctrl_inst1.g0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_idle_4_LC_4_20_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_idle_4_LC_4_20_5 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.counter_idle_4_LC_4_20_5 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_4_LC_4_20_5  (
            .in0(N__3936),
            .in1(N__3637),
            .in2(N__3570),
            .in3(N__3567),
            .lcout(\fsm_ctrl_inst1.counter_idleZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6138),
            .ce(),
            .sr(N__5822));
    defparam \fsm_ctrl_inst1.current_state_RNI31NH_0_LC_4_20_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.current_state_RNI31NH_0_LC_4_20_6 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.current_state_RNI31NH_0_LC_4_20_6 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \fsm_ctrl_inst1.current_state_RNI31NH_0_LC_4_20_6  (
            .in0(N__4690),
            .in1(N__4541),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fsm_ctrl_inst1.current_state_20_d_i ),
            .ltout(\fsm_ctrl_inst1.current_state_20_d_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_idle_2_LC_4_20_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_idle_2_LC_4_20_7 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.counter_idle_2_LC_4_20_7 .LUT_INIT=16'b1000111110001000;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_2_LC_4_20_7  (
            .in0(N__3561),
            .in1(N__3555),
            .in2(N__3549),
            .in3(N__3546),
            .lcout(\fsm_ctrl_inst1.counter_idleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6138),
            .ce(),
            .sr(N__5822));
    defparam \fsm_ctrl_inst1.current_state_RNO_0_0_LC_4_21_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.current_state_RNO_0_0_LC_4_21_0 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.current_state_RNO_0_0_LC_4_21_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fsm_ctrl_inst1.current_state_RNO_0_0_LC_4_21_0  (
            .in0(_gnd_net_),
            .in1(N__3968),
            .in2(_gnd_net_),
            .in3(N__4026),
            .lcout(),
            .ltout(\fsm_ctrl_inst1.N_93_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.current_state_0_LC_4_21_1 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.current_state_0_LC_4_21_1 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.current_state_0_LC_4_21_1 .LUT_INIT=16'b0001000100010000;
    LogicCell40 \fsm_ctrl_inst1.current_state_0_LC_4_21_1  (
            .in0(N__4852),
            .in1(N__3924),
            .in2(N__3540),
            .in3(N__4584),
            .lcout(fsm_ctrl_inst1_current_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6142),
            .ce(),
            .sr(N__5827));
    defparam \fsm_ctrl_inst1.counter_idle_RNO_1_0_LC_4_21_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_1_0_LC_4_21_4 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_1_0_LC_4_21_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_RNO_1_0_LC_4_21_4  (
            .in0(N__4076),
            .in1(N__3967),
            .in2(N__4014),
            .in3(N__4118),
            .lcout(),
            .ltout(\fsm_ctrl_inst1.counter_idle_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_idle_RNO_0_0_LC_4_21_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_0_0_LC_4_21_5 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_0_0_LC_4_21_5 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_RNO_0_0_LC_4_21_5  (
            .in0(_gnd_net_),
            .in1(N__4694),
            .in2(N__3666),
            .in3(N__4583),
            .lcout(),
            .ltout(\fsm_ctrl_inst1.counter_idlee_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_idle_0_LC_4_21_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_idle_0_LC_4_21_6 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.counter_idle_0_LC_4_21_6 .LUT_INIT=16'b1111000100000100;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_0_LC_4_21_6  (
            .in0(N__3639),
            .in1(N__3600),
            .in2(N__3663),
            .in3(N__4044),
            .lcout(\fsm_ctrl_inst1.counter_idleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6142),
            .ce(),
            .sr(N__5827));
    defparam \fsm_ctrl_inst1.counter_idle_1_LC_4_21_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_idle_1_LC_4_21_7 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.counter_idle_1_LC_4_21_7 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_1_LC_4_21_7  (
            .in0(N__3660),
            .in1(N__3654),
            .in2(N__3648),
            .in3(N__3638),
            .lcout(\fsm_ctrl_inst1.counter_idleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6142),
            .ce(),
            .sr(N__5827));
    defparam \fsm_ctrl_inst1.MOSI_LC_4_22_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.MOSI_LC_4_22_0 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.MOSI_LC_4_22_0 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \fsm_ctrl_inst1.MOSI_LC_4_22_0  (
            .in0(N__3621),
            .in1(N__4553),
            .in2(N__3615),
            .in3(N__4807),
            .lcout(MOSI),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6144),
            .ce(),
            .sr(N__5828));
    defparam CONSTANT_ONE_LUT4_LC_4_24_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_4_24_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_4_24_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_4_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_67_LC_5_13_1 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_67_LC_5_13_1 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_67_LC_5_13_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_67_LC_5_13_1  (
            .in0(N__5052),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3720),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6145),
            .ce(N__4217),
            .sr(N__5823));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_68_LC_5_13_2 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_68_LC_5_13_2 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_68_LC_5_13_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_68_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(N__3591),
            .in2(_gnd_net_),
            .in3(N__5053),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6145),
            .ce(N__4217),
            .sr(N__5823));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_65_LC_5_13_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_65_LC_5_13_3 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_65_LC_5_13_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_65_LC_5_13_3  (
            .in0(N__5050),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3585),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6145),
            .ce(N__4217),
            .sr(N__5823));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_64_LC_5_13_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_64_LC_5_13_6 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_64_LC_5_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_64_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(N__3753),
            .in2(_gnd_net_),
            .in3(N__5049),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6145),
            .ce(N__4217),
            .sr(N__5823));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_66_LC_5_13_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_66_LC_5_13_7 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_66_LC_5_13_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_66_LC_5_13_7  (
            .in0(N__5051),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3726),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6145),
            .ce(N__4217),
            .sr(N__5823));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_69_LC_5_14_1 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_69_LC_5_14_1 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_69_LC_5_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_69_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(N__3714),
            .in2(_gnd_net_),
            .in3(N__5045),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6143),
            .ce(N__4216),
            .sr(N__5818));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_70_LC_5_14_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_70_LC_5_14_5 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_70_LC_5_14_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_70_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(N__3708),
            .in2(_gnd_net_),
            .in3(N__5046),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6143),
            .ce(N__4216),
            .sr(N__5818));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_71_LC_5_14_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_71_LC_5_14_6 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_71_LC_5_14_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_71_LC_5_14_6  (
            .in0(N__5047),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3702),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6143),
            .ce(N__4216),
            .sr(N__5818));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_73_LC_5_15_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_73_LC_5_15_0 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_73_LC_5_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_73_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(N__3678),
            .in2(_gnd_net_),
            .in3(N__5008),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6139),
            .ce(N__4214),
            .sr(N__5814));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_74_LC_5_15_1 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_74_LC_5_15_1 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_74_LC_5_15_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_74_LC_5_15_1  (
            .in0(N__5009),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3696),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6139),
            .ce(N__4214),
            .sr(N__5814));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_19_LC_5_15_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_19_LC_5_15_4 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_19_LC_5_15_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_19_LC_5_15_4  (
            .in0(_gnd_net_),
            .in1(N__3672),
            .in2(_gnd_net_),
            .in3(N__5006),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6139),
            .ce(N__4214),
            .sr(N__5814));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_72_LC_5_15_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_72_LC_5_15_5 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_72_LC_5_15_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_72_LC_5_15_5  (
            .in0(N__5007),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3684),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6139),
            .ce(N__4214),
            .sr(N__5814));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_18_LC_5_15_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_18_LC_5_15_6 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_18_LC_5_15_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_18_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(N__3783),
            .in2(_gnd_net_),
            .in3(N__5005),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6139),
            .ce(N__4214),
            .sr(N__5814));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_14_LC_5_16_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_14_LC_5_16_0 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_14_LC_5_16_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_14_LC_5_16_0  (
            .in0(_gnd_net_),
            .in1(N__3831),
            .in2(_gnd_net_),
            .in3(N__4993),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6134),
            .ce(N__4212),
            .sr(N__5806));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_17_LC_5_16_1 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_17_LC_5_16_1 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_17_LC_5_16_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_17_LC_5_16_1  (
            .in0(N__4996),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3777),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6134),
            .ce(N__4212),
            .sr(N__5806));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_16_LC_5_16_2 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_16_LC_5_16_2 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_16_LC_5_16_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_16_LC_5_16_2  (
            .in0(_gnd_net_),
            .in1(N__3765),
            .in2(_gnd_net_),
            .in3(N__4995),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6134),
            .ce(N__4212),
            .sr(N__5806));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_21_LC_5_16_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_21_LC_5_16_3 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_21_LC_5_16_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_21_LC_5_16_3  (
            .in0(N__4997),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4227),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6134),
            .ce(N__4212),
            .sr(N__5806));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_15_LC_5_16_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_15_LC_5_16_5 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_15_LC_5_16_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_15_LC_5_16_5  (
            .in0(N__4994),
            .in1(N__3771),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6134),
            .ce(N__4212),
            .sr(N__5806));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_63_LC_5_16_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_63_LC_5_16_6 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_63_LC_5_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_63_LC_5_16_6  (
            .in0(_gnd_net_),
            .in1(N__3759),
            .in2(_gnd_net_),
            .in3(N__4999),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6134),
            .ce(N__4212),
            .sr(N__5806));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_22_LC_5_16_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_22_LC_5_16_7 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_22_LC_5_16_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_22_LC_5_16_7  (
            .in0(N__4998),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3744),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6134),
            .ce(N__4212),
            .sr(N__5806));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_27_LC_5_17_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_27_LC_5_17_0 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_27_LC_5_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_27_LC_5_17_0  (
            .in0(_gnd_net_),
            .in1(N__3846),
            .in2(_gnd_net_),
            .in3(N__4953),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6126),
            .ce(N__4205),
            .sr(N__5815));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_23_LC_5_17_1 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_23_LC_5_17_1 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_23_LC_5_17_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_23_LC_5_17_1  (
            .in0(N__4951),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3738),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6126),
            .ce(N__4205),
            .sr(N__5815));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_49_LC_5_17_2 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_49_LC_5_17_2 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_49_LC_5_17_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_49_LC_5_17_2  (
            .in0(_gnd_net_),
            .in1(N__3732),
            .in2(_gnd_net_),
            .in3(N__4954),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6126),
            .ce(N__4205),
            .sr(N__5815));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_26_LC_5_17_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_26_LC_5_17_3 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_26_LC_5_17_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_26_LC_5_17_3  (
            .in0(N__4952),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3807),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6126),
            .ce(N__4205),
            .sr(N__5815));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_13_LC_5_17_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_13_LC_5_17_4 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_13_LC_5_17_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_13_LC_5_17_4  (
            .in0(_gnd_net_),
            .in1(N__3840),
            .in2(_gnd_net_),
            .in3(N__4950),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6126),
            .ce(N__4205),
            .sr(N__5815));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_50_LC_5_17_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_50_LC_5_17_6 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_50_LC_5_17_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_50_LC_5_17_6  (
            .in0(_gnd_net_),
            .in1(N__3825),
            .in2(_gnd_net_),
            .in3(N__4955),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6126),
            .ce(N__4205),
            .sr(N__5815));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_51_LC_5_17_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_51_LC_5_17_7 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_51_LC_5_17_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_51_LC_5_17_7  (
            .in0(N__4956),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3819),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6126),
            .ce(N__4205),
            .sr(N__5815));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_47_LC_5_18_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_47_LC_5_18_0 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_47_LC_5_18_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_47_LC_5_18_0  (
            .in0(N__4948),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3900),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6135),
            .ce(N__4213),
            .sr(N__5819));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_25_LC_5_18_1 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_25_LC_5_18_1 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_25_LC_5_18_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_25_LC_5_18_1  (
            .in0(_gnd_net_),
            .in1(N__3912),
            .in2(_gnd_net_),
            .in3(N__4943),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6135),
            .ce(N__4213),
            .sr(N__5819));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_45_LC_5_18_2 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_45_LC_5_18_2 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_45_LC_5_18_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_45_LC_5_18_2  (
            .in0(N__4946),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3801),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6135),
            .ce(N__4213),
            .sr(N__5819));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_29_LC_5_18_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_29_LC_5_18_3 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_29_LC_5_18_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_29_LC_5_18_3  (
            .in0(_gnd_net_),
            .in1(N__3888),
            .in2(_gnd_net_),
            .in3(N__4945),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6135),
            .ce(N__4213),
            .sr(N__5819));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_52_LC_5_18_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_52_LC_5_18_4 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_52_LC_5_18_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_52_LC_5_18_4  (
            .in0(N__4949),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3795),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6135),
            .ce(N__4213),
            .sr(N__5819));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_24_LC_5_18_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_24_LC_5_18_5 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_24_LC_5_18_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_24_LC_5_18_5  (
            .in0(_gnd_net_),
            .in1(N__3918),
            .in2(_gnd_net_),
            .in3(N__4942),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6135),
            .ce(N__4213),
            .sr(N__5819));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_46_LC_5_18_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_46_LC_5_18_6 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_46_LC_5_18_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_46_LC_5_18_6  (
            .in0(N__4947),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3906),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6135),
            .ce(N__4213),
            .sr(N__5819));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_28_LC_5_18_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_28_LC_5_18_7 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_28_LC_5_18_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_28_LC_5_18_7  (
            .in0(_gnd_net_),
            .in1(N__3894),
            .in2(_gnd_net_),
            .in3(N__4944),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6135),
            .ce(N__4213),
            .sr(N__5819));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_33_LC_5_19_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_33_LC_5_19_0 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_33_LC_5_19_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_33_LC_5_19_0  (
            .in0(_gnd_net_),
            .in1(N__4128),
            .in2(_gnd_net_),
            .in3(N__4864),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6140),
            .ce(N__4215),
            .sr(N__5824));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_34_LC_5_19_1 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_34_LC_5_19_1 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_34_LC_5_19_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_34_LC_5_19_1  (
            .in0(N__4865),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3882),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6140),
            .ce(N__4215),
            .sr(N__5824));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_30_LC_5_19_2 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_30_LC_5_19_2 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_30_LC_5_19_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_30_LC_5_19_2  (
            .in0(_gnd_net_),
            .in1(N__3876),
            .in2(_gnd_net_),
            .in3(N__4861),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6140),
            .ce(N__4215),
            .sr(N__5824));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_35_LC_5_19_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_35_LC_5_19_3 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_35_LC_5_19_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_35_LC_5_19_3  (
            .in0(N__4866),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3870),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6140),
            .ce(N__4215),
            .sr(N__5824));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_31_LC_5_19_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_31_LC_5_19_5 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_31_LC_5_19_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_31_LC_5_19_5  (
            .in0(N__4862),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3864),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6140),
            .ce(N__4215),
            .sr(N__5824));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_36_LC_5_19_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_36_LC_5_19_6 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_36_LC_5_19_6 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_36_LC_5_19_6  (
            .in0(_gnd_net_),
            .in1(N__3858),
            .in2(_gnd_net_),
            .in3(N__4867),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6140),
            .ce(N__4215),
            .sr(N__5824));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_32_LC_5_19_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_32_LC_5_19_7 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_32_LC_5_19_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_32_LC_5_19_7  (
            .in0(N__4863),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4134),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6140),
            .ce(N__4215),
            .sr(N__5824));
    defparam \fsm_ctrl_inst1.current_state_RNO_2_0_LC_5_20_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.current_state_RNO_2_0_LC_5_20_0 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.current_state_RNO_2_0_LC_5_20_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \fsm_ctrl_inst1.current_state_RNO_2_0_LC_5_20_0  (
            .in0(N__4117),
            .in1(N__4074),
            .in2(N__4013),
            .in3(N__4043),
            .lcout(\fsm_ctrl_inst1.current_state_RNO_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_idle_RNO_2_3_LC_5_20_2 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_2_3_LC_5_20_2 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_2_3_LC_5_20_2 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_RNO_2_3_LC_5_20_2  (
            .in0(N__4005),
            .in1(N__3970),
            .in2(N__4809),
            .in3(N__4508),
            .lcout(\fsm_ctrl_inst1.g0_0_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \config_register_latched_dec_inst1.STATSR_cnv_x0_0_LC_5_20_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_cnv_x0_0_LC_5_20_4 .SEQ_MODE=4'b0000;
    defparam \config_register_latched_dec_inst1.STATSR_cnv_x0_0_LC_5_20_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_cnv_x0_0_LC_5_20_4  (
            .in0(N__5093),
            .in1(N__4439),
            .in2(N__5076),
            .in3(N__4507),
            .lcout(\config_register_latched_dec_inst1.STATSR_cnv_x0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_idle_RNO_2_4_LC_5_20_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_2_4_LC_5_20_6 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.counter_idle_RNO_2_4_LC_5_20_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \fsm_ctrl_inst1.counter_idle_RNO_2_4_LC_5_20_6  (
            .in0(N__4006),
            .in1(N__3971),
            .in2(N__4810),
            .in3(N__4509),
            .lcout(\fsm_ctrl_inst1.g0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_din_RNO_0_3_LC_5_21_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_din_RNO_0_3_LC_5_21_0 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.counter_din_RNO_0_3_LC_5_21_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \fsm_ctrl_inst1.counter_din_RNO_0_3_LC_5_21_0  (
            .in0(N__4327),
            .in1(N__4272),
            .in2(N__4313),
            .in3(N__4287),
            .lcout(),
            .ltout(\fsm_ctrl_inst1.counter_din_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_din_3_LC_5_21_1 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_din_3_LC_5_21_1 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.counter_din_3_LC_5_21_1 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \fsm_ctrl_inst1.counter_din_3_LC_5_21_1  (
            .in0(N__4567),
            .in1(_gnd_net_),
            .in2(N__3930),
            .in3(_gnd_net_),
            .lcout(\fsm_ctrl_inst1.counter_dinZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6146),
            .ce(),
            .sr(N__5829));
    defparam \fsm_ctrl_inst1.current_state_RNO_3_0_LC_5_21_2 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.current_state_RNO_3_0_LC_5_21_2 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.current_state_RNO_3_0_LC_5_21_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \fsm_ctrl_inst1.current_state_RNO_3_0_LC_5_21_2  (
            .in0(N__4326),
            .in1(N__4565),
            .in2(N__4312),
            .in3(N__4286),
            .lcout(),
            .ltout(\fsm_ctrl_inst1.current_state_RNO_3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.current_state_RNO_1_0_LC_5_21_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.current_state_RNO_1_0_LC_5_21_3 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.current_state_RNO_1_0_LC_5_21_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \fsm_ctrl_inst1.current_state_RNO_1_0_LC_5_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3927),
            .in3(N__4268),
            .lcout(\fsm_ctrl_inst1.current_state_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.counter_din_1_LC_5_21_4 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_din_1_LC_5_21_4 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.counter_din_1_LC_5_21_4 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \fsm_ctrl_inst1.counter_din_1_LC_5_21_4  (
            .in0(N__4269),
            .in1(N__4569),
            .in2(_gnd_net_),
            .in3(N__4288),
            .lcout(\fsm_ctrl_inst1.counter_dinZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6146),
            .ce(),
            .sr(N__5829));
    defparam \fsm_ctrl_inst1.counter_din_2_LC_5_21_5 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.counter_din_2_LC_5_21_5 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.counter_din_2_LC_5_21_5 .LUT_INIT=16'b0010101010000000;
    LogicCell40 \fsm_ctrl_inst1.counter_din_2_LC_5_21_5  (
            .in0(N__4568),
            .in1(N__4270),
            .in2(N__4293),
            .in3(N__4329),
            .lcout(\fsm_ctrl_inst1.counter_dinZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6146),
            .ce(),
            .sr(N__5829));
    defparam \fsm_ctrl_inst1.current_state_RNO_0_1_LC_5_21_6 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.current_state_RNO_0_1_LC_5_21_6 .SEQ_MODE=4'b0000;
    defparam \fsm_ctrl_inst1.current_state_RNO_0_1_LC_5_21_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \fsm_ctrl_inst1.current_state_RNO_0_1_LC_5_21_6  (
            .in0(N__4328),
            .in1(_gnd_net_),
            .in2(N__4314),
            .in3(N__4566),
            .lcout(),
            .ltout(\fsm_ctrl_inst1.o2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.current_state_1_LC_5_21_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.current_state_1_LC_5_21_7 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.current_state_1_LC_5_21_7 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \fsm_ctrl_inst1.current_state_1_LC_5_21_7  (
            .in0(N__4292),
            .in1(N__4271),
            .in2(N__4242),
            .in3(N__4806),
            .lcout(fsm_ctrl_inst1_current_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6146),
            .ce(),
            .sr(N__5829));
    defparam \config_register_latched_dec_inst1.STATSR_0_LC_5_23_1 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_0_LC_5_23_1 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_0_LC_5_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_0_LC_5_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4418),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6150),
            .ce(N__5976),
            .sr(N__5832));
    defparam \config_register_latched_dec_inst1.STATSR_1_LC_5_24_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_1_LC_5_24_6 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_1_LC_5_24_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_1_LC_5_24_6  (
            .in0(_gnd_net_),
            .in1(N__4239),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6153),
            .ce(N__5975),
            .sr(N__5835));
    defparam \fsm_ctrl_inst1.bit_sequence_stat_20_LC_6_14_0 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_20_LC_6_14_0 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.bit_sequence_stat_20_LC_6_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fsm_ctrl_inst1.bit_sequence_stat_20_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(N__4233),
            .in2(_gnd_net_),
            .in3(N__5048),
            .lcout(\fsm_ctrl_inst1.bit_sequence_statZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6147),
            .ce(N__4218),
            .sr(N__5825));
    defparam \config_register_latched_dec_inst1.DYNSR_RNIQ2U9_15_LC_6_19_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_RNIQ2U9_15_LC_6_19_6 .SEQ_MODE=4'b0000;
    defparam \config_register_latched_dec_inst1.DYNSR_RNIQ2U9_15_LC_6_19_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_RNIQ2U9_15_LC_6_19_6  (
            .in0(N__4368),
            .in1(N__5202),
            .in2(_gnd_net_),
            .in3(N__4446),
            .lcout(SDO_signal_out_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \config_register_latched_dec_inst1.DYNSR_12_LC_6_20_0 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_12_LC_6_20_0 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.DYNSR_12_LC_6_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_12_LC_6_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4344),
            .lcout(\config_register_latched_dec_inst1.DYNSRZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6148),
            .ce(N__5145),
            .sr(N__5830));
    defparam \config_register_latched_dec_inst1.DYNSR_14_LC_6_20_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_14_LC_6_20_3 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.DYNSR_14_LC_6_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_14_LC_6_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4356),
            .lcout(\config_register_latched_dec_inst1.DYNSRZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6148),
            .ce(N__5145),
            .sr(N__5830));
    defparam \config_register_latched_dec_inst1.DYNSR_10_LC_6_20_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_10_LC_6_20_4 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.DYNSR_10_LC_6_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_10_LC_6_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5193),
            .lcout(\config_register_latched_dec_inst1.DYNSRZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6148),
            .ce(N__5145),
            .sr(N__5830));
    defparam \config_register_latched_dec_inst1.DYNSR_15_LC_6_20_5 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_15_LC_6_20_5 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.DYNSR_15_LC_6_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_15_LC_6_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4374),
            .lcout(\config_register_latched_dec_inst1.DYNSRZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6148),
            .ce(N__5145),
            .sr(N__5830));
    defparam \config_register_latched_dec_inst1.DYNSR_13_LC_6_20_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_13_LC_6_20_6 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.DYNSR_13_LC_6_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_13_LC_6_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4362),
            .lcout(\config_register_latched_dec_inst1.DYNSRZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6148),
            .ce(N__5145),
            .sr(N__5830));
    defparam \config_register_latched_dec_inst1.DYNSR_11_LC_6_20_7 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_11_LC_6_20_7 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.DYNSR_11_LC_6_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_11_LC_6_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4350),
            .lcout(\config_register_latched_dec_inst1.DYNSRZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6148),
            .ce(N__5145),
            .sr(N__5830));
    defparam \config_register_latched_dec_inst1.DYNSR_cnv_x0_0_LC_6_21_0 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_cnv_x0_0_LC_6_21_0 .SEQ_MODE=4'b0000;
    defparam \config_register_latched_dec_inst1.DYNSR_cnv_x0_0_LC_6_21_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_cnv_x0_0_LC_6_21_0  (
            .in0(N__4554),
            .in1(N__5075),
            .in2(N__5115),
            .in3(N__4442),
            .lcout(),
            .ltout(\config_register_latched_dec_inst1.DYNSR_cnv_x0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \config_register_latched_dec_inst1.DYNSR_cnv_ns_0_LC_6_21_1 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_cnv_ns_0_LC_6_21_1 .SEQ_MODE=4'b0000;
    defparam \config_register_latched_dec_inst1.DYNSR_cnv_ns_0_LC_6_21_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_cnv_ns_0_LC_6_21_1  (
            .in0(_gnd_net_),
            .in1(N__4335),
            .in2(N__4338),
            .in3(N__4688),
            .lcout(\config_register_latched_dec_inst1.DYNSR_cnv_nsZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \config_register_latched_dec_inst1.DYNSR_cnv_x1_0_LC_6_21_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_cnv_x1_0_LC_6_21_2 .SEQ_MODE=4'b0000;
    defparam \config_register_latched_dec_inst1.DYNSR_cnv_x1_0_LC_6_21_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_cnv_x1_0_LC_6_21_2  (
            .in0(N__5112),
            .in1(N__5073),
            .in2(_gnd_net_),
            .in3(N__4440),
            .lcout(\config_register_latched_dec_inst1.DYNSR_cnv_x1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.SCLK_LC_6_21_3 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.SCLK_LC_6_21_3 .SEQ_MODE=4'b1010;
    defparam \fsm_ctrl_inst1.SCLK_LC_6_21_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \fsm_ctrl_inst1.SCLK_LC_6_21_3  (
            .in0(N__5114),
            .in1(N__4689),
            .in2(_gnd_net_),
            .in3(N__4556),
            .lcout(fsm_ctrl_inst1_SCLK_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6149),
            .ce(),
            .sr(N__5831));
    defparam \config_register_latched_dec_inst1.STATSR_cnv_x1_0_LC_6_21_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_cnv_x1_0_LC_6_21_4 .SEQ_MODE=4'b0000;
    defparam \config_register_latched_dec_inst1.STATSR_cnv_x1_0_LC_6_21_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_cnv_x1_0_LC_6_21_4  (
            .in0(N__5113),
            .in1(N__4441),
            .in2(_gnd_net_),
            .in3(N__5074),
            .lcout(),
            .ltout(\config_register_latched_dec_inst1.STATSR_cnv_x1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \config_register_latched_dec_inst1.STATSR_cnv_ns_0_LC_6_21_5 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_cnv_ns_0_LC_6_21_5 .SEQ_MODE=4'b0000;
    defparam \config_register_latched_dec_inst1.STATSR_cnv_ns_0_LC_6_21_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_cnv_ns_0_LC_6_21_5  (
            .in0(_gnd_net_),
            .in1(N__4687),
            .in2(N__4617),
            .in3(N__4614),
            .lcout(STATSR_cnv_ns_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fsm_ctrl_inst1.SEL_LC_6_21_7 .C_ON=1'b0;
    defparam \fsm_ctrl_inst1.SEL_LC_6_21_7 .SEQ_MODE=4'b1011;
    defparam \fsm_ctrl_inst1.SEL_LC_6_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \fsm_ctrl_inst1.SEL_LC_6_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4555),
            .lcout(SEL_REG),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6149),
            .ce(),
            .sr(N__5831));
    defparam \config_register_latched_dec_inst1.DYNSR_2_LC_6_22_0 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_2_LC_6_22_0 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.DYNSR_2_LC_6_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_2_LC_6_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4398),
            .lcout(\config_register_latched_dec_inst1.DYNSRZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6151),
            .ce(N__5153),
            .sr(N__5833));
    defparam \config_register_latched_dec_inst1.DYNSR_0_LC_6_22_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_0_LC_6_22_4 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.DYNSR_0_LC_6_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_0_LC_6_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4419),
            .lcout(\config_register_latched_dec_inst1.DYNSRZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6151),
            .ce(N__5153),
            .sr(N__5833));
    defparam \config_register_latched_dec_inst1.DYNSR_1_LC_6_22_5 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_1_LC_6_22_5 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.DYNSR_1_LC_6_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_1_LC_6_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4404),
            .lcout(\config_register_latched_dec_inst1.DYNSRZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6151),
            .ce(N__5153),
            .sr(N__5833));
    defparam \config_register_latched_dec_inst1.DYNSR_3_LC_6_22_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_3_LC_6_22_6 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.DYNSR_3_LC_6_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_3_LC_6_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4392),
            .lcout(\config_register_latched_dec_inst1.DYNSRZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6151),
            .ce(N__5153),
            .sr(N__5833));
    defparam \config_register_latched_dec_inst1.DYNSR_4_LC_6_22_7 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_4_LC_6_22_7 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.DYNSR_4_LC_6_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_4_LC_6_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4386),
            .lcout(\config_register_latched_dec_inst1.DYNSRZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6151),
            .ce(N__5153),
            .sr(N__5833));
    defparam \config_register_latched_dec_inst1.STATSR_2_LC_6_24_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_2_LC_6_24_3 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_2_LC_6_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_2_LC_6_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4380),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6155),
            .ce(N__5974),
            .sr(N__5837));
    defparam \config_register_latched_dec_inst1.STATSR_3_LC_6_24_5 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_3_LC_6_24_5 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_3_LC_6_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_3_LC_6_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5214),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6155),
            .ce(N__5974),
            .sr(N__5837));
    defparam \config_register_latched_dec_inst1.STATSR_4_LC_6_24_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_4_LC_6_24_6 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_4_LC_6_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_4_LC_6_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5208),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6155),
            .ce(N__5974),
            .sr(N__5837));
    defparam \config_register_latched_dec_inst1.STATSR_87_LC_6_25_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_87_LC_6_25_2 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_87_LC_6_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_87_LC_6_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5262),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6156),
            .ce(N__5972),
            .sr(N__5838));
    defparam \config_register_latched_dec_inst1.DYNSR_9_LC_7_21_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_9_LC_7_21_2 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.DYNSR_9_LC_7_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_9_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5175),
            .lcout(\config_register_latched_dec_inst1.DYNSRZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6152),
            .ce(N__5157),
            .sr(N__5834));
    defparam \config_register_latched_dec_inst1.DYNSR_6_LC_7_21_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_6_LC_7_21_3 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.DYNSR_6_LC_7_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_6_LC_7_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5163),
            .lcout(\config_register_latched_dec_inst1.DYNSRZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6152),
            .ce(N__5157),
            .sr(N__5834));
    defparam \config_register_latched_dec_inst1.DYNSR_7_LC_7_21_5 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_7_LC_7_21_5 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.DYNSR_7_LC_7_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_7_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5187),
            .lcout(\config_register_latched_dec_inst1.DYNSRZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6152),
            .ce(N__5157),
            .sr(N__5834));
    defparam \config_register_latched_dec_inst1.DYNSR_8_LC_7_21_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_8_LC_7_21_6 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.DYNSR_8_LC_7_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_8_LC_7_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5181),
            .lcout(\config_register_latched_dec_inst1.DYNSRZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6152),
            .ce(N__5157),
            .sr(N__5834));
    defparam \config_register_latched_dec_inst1.DYNSR_5_LC_7_22_5 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.DYNSR_5_LC_7_22_5 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.DYNSR_5_LC_7_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.DYNSR_5_LC_7_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5169),
            .lcout(\config_register_latched_dec_inst1.DYNSRZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6154),
            .ce(N__5152),
            .sr(N__5836));
    defparam \config_register_latched_dec_inst1.STATSR_6_LC_7_24_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_6_LC_7_24_2 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_6_LC_7_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_6_LC_7_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5268),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6157),
            .ce(N__5973),
            .sr(N__5839));
    defparam \config_register_latched_dec_inst1.STATSR_5_LC_7_24_7 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_5_LC_7_24_7 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_5_LC_7_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_5_LC_7_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5274),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6157),
            .ce(N__5973),
            .sr(N__5839));
    defparam \config_register_latched_dec_inst1.STATSR_86_LC_7_25_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_86_LC_7_25_6 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_86_LC_7_25_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_86_LC_7_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5229),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6158),
            .ce(N__5971),
            .sr(N__5840));
    defparam \config_register_latched_dec_inst1.STATSR_8_LC_9_24_0 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_8_LC_9_24_0 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_8_LC_9_24_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_8_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5247),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6159),
            .ce(N__5970),
            .sr(N__5841));
    defparam \config_register_latched_dec_inst1.STATSR_7_LC_9_24_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_7_LC_9_24_4 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_7_LC_9_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_7_LC_9_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5256),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6159),
            .ce(N__5970),
            .sr(N__5841));
    defparam \config_register_latched_dec_inst1.STATSR_84_LC_9_25_0 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_84_LC_9_25_0 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_84_LC_9_25_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_84_LC_9_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5316),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6160),
            .ce(N__5969),
            .sr(N__5842));
    defparam \config_register_latched_dec_inst1.STATSR_9_LC_9_25_1 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_9_LC_9_25_1 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_9_LC_9_25_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_9_LC_9_25_1  (
            .in0(_gnd_net_),
            .in1(N__5241),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6160),
            .ce(N__5969),
            .sr(N__5842));
    defparam \config_register_latched_dec_inst1.STATSR_85_LC_9_25_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_85_LC_9_25_3 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_85_LC_9_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_85_LC_9_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5235),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6160),
            .ce(N__5969),
            .sr(N__5842));
    defparam \config_register_latched_dec_inst1.STATSR_12_LC_10_25_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_12_LC_10_25_3 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_12_LC_10_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_12_LC_10_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5322),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6161),
            .ce(N__5968),
            .sr(N__5843));
    defparam \config_register_latched_dec_inst1.STATSR_10_LC_10_25_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_10_LC_10_25_4 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_10_LC_10_25_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_10_LC_10_25_4  (
            .in0(_gnd_net_),
            .in1(N__5220),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6161),
            .ce(N__5968),
            .sr(N__5843));
    defparam \config_register_latched_dec_inst1.STATSR_11_LC_10_25_7 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_11_LC_10_25_7 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_11_LC_10_25_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_11_LC_10_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5328),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6161),
            .ce(N__5968),
            .sr(N__5843));
    defparam \config_register_latched_dec_inst1.STATSR_83_LC_10_26_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_83_LC_10_26_6 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_83_LC_10_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_83_LC_10_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5298),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6162),
            .ce(N__5966),
            .sr(N__5844));
    defparam \config_register_latched_dec_inst1.STATSR_13_LC_11_25_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_13_LC_11_25_2 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_13_LC_11_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_13_LC_11_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5310),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6163),
            .ce(N__5967),
            .sr(N__5845));
    defparam \config_register_latched_dec_inst1.STATSR_81_LC_11_26_5 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_81_LC_11_26_5 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_81_LC_11_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_81_LC_11_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5286),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6164),
            .ce(N__5964),
            .sr(N__5846));
    defparam \config_register_latched_dec_inst1.STATSR_82_LC_11_26_7 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_82_LC_11_26_7 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_82_LC_11_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_82_LC_11_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5304),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6164),
            .ce(N__5964),
            .sr(N__5846));
    defparam \config_register_latched_dec_inst1.STATSR_14_LC_12_25_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_14_LC_12_25_2 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_14_LC_12_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_14_LC_12_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5292),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6165),
            .ce(N__5965),
            .sr(N__5847));
    defparam \config_register_latched_dec_inst1.STATSR_77_LC_12_27_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_77_LC_12_27_2 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_77_LC_12_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_77_LC_12_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5364),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6167),
            .ce(N__5961),
            .sr(N__5849));
    defparam \config_register_latched_dec_inst1.STATSR_80_LC_12_27_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_80_LC_12_27_3 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_80_LC_12_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_80_LC_12_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5280),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6167),
            .ce(N__5961),
            .sr(N__5849));
    defparam \config_register_latched_dec_inst1.STATSR_79_LC_12_27_5 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_79_LC_12_27_5 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_79_LC_12_27_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_79_LC_12_27_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5382),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6167),
            .ce(N__5961),
            .sr(N__5849));
    defparam \config_register_latched_dec_inst1.STATSR_78_LC_12_27_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_78_LC_12_27_6 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_78_LC_12_27_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_78_LC_12_27_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5388),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6167),
            .ce(N__5961),
            .sr(N__5849));
    defparam \config_register_latched_dec_inst1.STATSR_15_LC_13_25_1 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_15_LC_13_25_1 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_15_LC_13_25_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_15_LC_13_25_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5376),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6166),
            .ce(N__5963),
            .sr(N__5848));
    defparam \config_register_latched_dec_inst1.STATSR_75_LC_13_27_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_75_LC_13_27_2 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_75_LC_13_27_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_75_LC_13_27_2  (
            .in0(_gnd_net_),
            .in1(N__5358),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6169),
            .ce(N__5959),
            .sr(N__5851));
    defparam \config_register_latched_dec_inst1.STATSR_76_LC_13_27_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_76_LC_13_27_3 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_76_LC_13_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_76_LC_13_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5370),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6169),
            .ce(N__5959),
            .sr(N__5851));
    defparam \config_register_latched_dec_inst1.STATSR_74_LC_13_28_1 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_74_LC_13_28_1 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_74_LC_13_28_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_74_LC_13_28_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5340),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6171),
            .ce(N__5957),
            .sr(N__5853));
    defparam \config_register_latched_dec_inst1.STATSR_16_LC_14_25_1 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_16_LC_14_25_1 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_16_LC_14_25_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_16_LC_14_25_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5352),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6168),
            .ce(N__5962),
            .sr(N__5850));
    defparam \config_register_latched_dec_inst1.STATSR_17_LC_14_26_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_17_LC_14_26_3 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_17_LC_14_26_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_17_LC_14_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5346),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6170),
            .ce(N__5960),
            .sr(N__5852));
    defparam \config_register_latched_dec_inst1.STATSR_73_LC_14_28_1 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_73_LC_14_28_1 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_73_LC_14_28_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_73_LC_14_28_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5424),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6173),
            .ce(N__5956),
            .sr(N__5855));
    defparam \config_register_latched_dec_inst1.STATSR_18_LC_15_26_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_18_LC_15_26_2 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_18_LC_15_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_18_LC_15_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5334),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6172),
            .ce(N__5958),
            .sr(N__5854));
    defparam \config_register_latched_dec_inst1.STATSR_19_LC_15_26_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_19_LC_15_26_6 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_19_LC_15_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_19_LC_15_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5436),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6172),
            .ce(N__5958),
            .sr(N__5854));
    defparam \config_register_latched_dec_inst1.STATSR_71_LC_15_28_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_71_LC_15_28_2 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_71_LC_15_28_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_71_LC_15_28_2  (
            .in0(_gnd_net_),
            .in1(N__5418),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6174),
            .ce(N__5953),
            .sr(N__5856));
    defparam \config_register_latched_dec_inst1.STATSR_72_LC_15_28_5 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_72_LC_15_28_5 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_72_LC_15_28_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_72_LC_15_28_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5430),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6174),
            .ce(N__5953),
            .sr(N__5856));
    defparam \config_register_latched_dec_inst1.STATSR_70_LC_15_29_1 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_70_LC_15_29_1 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_70_LC_15_29_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_70_LC_15_29_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5406),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6176),
            .ce(N__5950),
            .sr(N__5858));
    defparam \config_register_latched_dec_inst1.STATSR_68_LC_15_29_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_68_LC_15_29_2 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_68_LC_15_29_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_68_LC_15_29_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5400),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6176),
            .ce(N__5950),
            .sr(N__5858));
    defparam \config_register_latched_dec_inst1.STATSR_69_LC_15_29_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_69_LC_15_29_3 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_69_LC_15_29_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_69_LC_15_29_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5412),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6176),
            .ce(N__5950),
            .sr(N__5858));
    defparam \config_register_latched_dec_inst1.STATSR_67_LC_15_29_7 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_67_LC_15_29_7 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_67_LC_15_29_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_67_LC_15_29_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5394),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6176),
            .ce(N__5950),
            .sr(N__5858));
    defparam \config_register_latched_dec_inst1.STATSR_66_LC_15_30_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_66_LC_15_30_4 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_66_LC_15_30_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_66_LC_15_30_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5442),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6179),
            .ce(N__5948),
            .sr(N__5861));
    defparam \config_register_latched_dec_inst1.STATSR_21_LC_16_27_0 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_21_LC_16_27_0 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_21_LC_16_27_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_21_LC_16_27_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5490),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6175),
            .ce(N__5954),
            .sr(N__5857));
    defparam \config_register_latched_dec_inst1.STATSR_20_LC_16_27_1 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_20_LC_16_27_1 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_20_LC_16_27_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_20_LC_16_27_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5496),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6175),
            .ce(N__5954),
            .sr(N__5857));
    defparam \config_register_latched_dec_inst1.STATSR_41_LC_16_27_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_41_LC_16_27_2 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_41_LC_16_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_41_LC_16_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5478),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6175),
            .ce(N__5954),
            .sr(N__5857));
    defparam \config_register_latched_dec_inst1.STATSR_42_LC_16_27_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_42_LC_16_27_3 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_42_LC_16_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_42_LC_16_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5484),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6175),
            .ce(N__5954),
            .sr(N__5857));
    defparam \config_register_latched_dec_inst1.STATSR_40_LC_16_27_5 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_40_LC_16_27_5 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_40_LC_16_27_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_40_LC_16_27_5  (
            .in0(N__5526),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6175),
            .ce(N__5954),
            .sr(N__5857));
    defparam \config_register_latched_dec_inst1.STATSR_44_LC_16_28_0 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_44_LC_16_28_0 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_44_LC_16_28_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_44_LC_16_28_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5466),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6177),
            .ce(N__5951),
            .sr(N__5859));
    defparam \config_register_latched_dec_inst1.STATSR_43_LC_16_28_1 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_43_LC_16_28_1 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_43_LC_16_28_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_43_LC_16_28_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5472),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6177),
            .ce(N__5951),
            .sr(N__5859));
    defparam \config_register_latched_dec_inst1.STATSR_45_LC_16_28_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_45_LC_16_28_3 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_45_LC_16_28_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_45_LC_16_28_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5460),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6177),
            .ce(N__5951),
            .sr(N__5859));
    defparam \config_register_latched_dec_inst1.STATSR_46_LC_16_28_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_46_LC_16_28_4 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_46_LC_16_28_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_46_LC_16_28_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5454),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6177),
            .ce(N__5951),
            .sr(N__5859));
    defparam \config_register_latched_dec_inst1.STATSR_22_LC_16_28_7 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_22_LC_16_28_7 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_22_LC_16_28_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_22_LC_16_28_7  (
            .in0(_gnd_net_),
            .in1(N__5448),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6177),
            .ce(N__5951),
            .sr(N__5859));
    defparam \config_register_latched_dec_inst1.STATSR_65_LC_16_30_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_65_LC_16_30_2 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_65_LC_16_30_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_65_LC_16_30_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5568),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6182),
            .ce(N__5945),
            .sr(N__5864));
    defparam \config_register_latched_dec_inst1.STATSR_36_LC_17_27_0 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_36_LC_17_27_0 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_36_LC_17_27_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_36_LC_17_27_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5544),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6178),
            .ce(N__5949),
            .sr(N__5860));
    defparam \config_register_latched_dec_inst1.STATSR_37_LC_17_27_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_37_LC_17_27_2 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_37_LC_17_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_37_LC_17_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5550),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6178),
            .ce(N__5949),
            .sr(N__5860));
    defparam \config_register_latched_dec_inst1.STATSR_35_LC_17_27_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_35_LC_17_27_3 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_35_LC_17_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_35_LC_17_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5640),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6178),
            .ce(N__5949),
            .sr(N__5860));
    defparam \config_register_latched_dec_inst1.STATSR_38_LC_17_27_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_38_LC_17_27_4 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_38_LC_17_27_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_38_LC_17_27_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5538),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6178),
            .ce(N__5949),
            .sr(N__5860));
    defparam \config_register_latched_dec_inst1.STATSR_39_LC_17_27_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_39_LC_17_27_6 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_39_LC_17_27_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_39_LC_17_27_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5532),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6178),
            .ce(N__5949),
            .sr(N__5860));
    defparam \config_register_latched_dec_inst1.STATSR_47_LC_17_28_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_47_LC_17_28_2 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_47_LC_17_28_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_47_LC_17_28_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5520),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6180),
            .ce(N__5947),
            .sr(N__5862));
    defparam \config_register_latched_dec_inst1.STATSR_48_LC_17_28_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_48_LC_17_28_4 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_48_LC_17_28_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_48_LC_17_28_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5514),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6180),
            .ce(N__5947),
            .sr(N__5862));
    defparam \config_register_latched_dec_inst1.STATSR_23_LC_17_28_5 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_23_LC_17_28_5 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_23_LC_17_28_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_23_LC_17_28_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5508),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6180),
            .ce(N__5947),
            .sr(N__5862));
    defparam \config_register_latched_dec_inst1.STATSR_49_LC_17_28_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_49_LC_17_28_6 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_49_LC_17_28_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_49_LC_17_28_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5502),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6180),
            .ce(N__5947),
            .sr(N__5862));
    defparam \config_register_latched_dec_inst1.STATSR_24_LC_17_28_7 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_24_LC_17_28_7 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_24_LC_17_28_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_24_LC_17_28_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5598),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6180),
            .ce(N__5947),
            .sr(N__5862));
    defparam \config_register_latched_dec_inst1.STATSR_50_LC_17_29_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_50_LC_17_29_2 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_50_LC_17_29_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_50_LC_17_29_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5592),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6183),
            .ce(N__5944),
            .sr(N__5865));
    defparam \config_register_latched_dec_inst1.STATSR_52_LC_17_29_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_52_LC_17_29_3 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_52_LC_17_29_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_52_LC_17_29_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5574),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6183),
            .ce(N__5944),
            .sr(N__5865));
    defparam \config_register_latched_dec_inst1.STATSR_53_LC_17_29_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_53_LC_17_29_4 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_53_LC_17_29_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_53_LC_17_29_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5586),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6183),
            .ce(N__5944),
            .sr(N__5865));
    defparam \config_register_latched_dec_inst1.STATSR_51_LC_17_29_7 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_51_LC_17_29_7 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_51_LC_17_29_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_51_LC_17_29_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5580),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6183),
            .ce(N__5944),
            .sr(N__5865));
    defparam \config_register_latched_dec_inst1.STATSR_64_LC_17_30_0 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_64_LC_17_30_0 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_64_LC_17_30_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_64_LC_17_30_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5562),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6185),
            .ce(N__5943),
            .sr(N__5867));
    defparam \config_register_latched_dec_inst1.STATSR_63_LC_17_30_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_63_LC_17_30_4 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_63_LC_17_30_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_63_LC_17_30_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5652),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6185),
            .ce(N__5943),
            .sr(N__5867));
    defparam \config_register_latched_dec_inst1.STATSR_61_LC_17_30_5 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_61_LC_17_30_5 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_61_LC_17_30_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_61_LC_17_30_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6228),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6185),
            .ce(N__5943),
            .sr(N__5867));
    defparam \config_register_latched_dec_inst1.STATSR_54_LC_17_30_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_54_LC_17_30_6 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_54_LC_17_30_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_54_LC_17_30_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5556),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6185),
            .ce(N__5943),
            .sr(N__5867));
    defparam \config_register_latched_dec_inst1.STATSR_62_LC_17_30_7 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_62_LC_17_30_7 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_62_LC_17_30_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_62_LC_17_30_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5658),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6185),
            .ce(N__5943),
            .sr(N__5867));
    defparam \config_register_latched_dec_inst1.STATSR_31_LC_18_27_1 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_31_LC_18_27_1 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_31_LC_18_27_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_31_LC_18_27_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5646),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6181),
            .ce(N__5955),
            .sr(N__5863));
    defparam \config_register_latched_dec_inst1.STATSR_30_LC_18_27_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_30_LC_18_27_2 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_30_LC_18_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_30_LC_18_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6234),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6181),
            .ce(N__5955),
            .sr(N__5863));
    defparam \config_register_latched_dec_inst1.STATSR_34_LC_18_27_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_34_LC_18_27_4 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_34_LC_18_27_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_34_LC_18_27_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5622),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6181),
            .ce(N__5955),
            .sr(N__5863));
    defparam \config_register_latched_dec_inst1.STATSR_32_LC_18_27_5 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_32_LC_18_27_5 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_32_LC_18_27_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_32_LC_18_27_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5634),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6181),
            .ce(N__5955),
            .sr(N__5863));
    defparam \config_register_latched_dec_inst1.STATSR_33_LC_18_27_7 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_33_LC_18_27_7 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_33_LC_18_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_33_LC_18_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5628),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6181),
            .ce(N__5955),
            .sr(N__5863));
    defparam \config_register_latched_dec_inst1.STATSR_26_LC_18_28_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_26_LC_18_28_3 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_26_LC_18_28_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_26_LC_18_28_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5604),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6184),
            .ce(N__5952),
            .sr(N__5866));
    defparam \config_register_latched_dec_inst1.STATSR_27_LC_18_28_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_27_LC_18_28_4 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_27_LC_18_28_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_27_LC_18_28_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5616),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6184),
            .ce(N__5952),
            .sr(N__5866));
    defparam \config_register_latched_dec_inst1.STATSR_25_LC_18_28_5 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_25_LC_18_28_5 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_25_LC_18_28_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_25_LC_18_28_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5610),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6184),
            .ce(N__5952),
            .sr(N__5866));
    defparam \config_register_latched_dec_inst1.STATSR_28_LC_18_28_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_28_LC_18_28_6 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_28_LC_18_28_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_28_LC_18_28_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6246),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6184),
            .ce(N__5952),
            .sr(N__5866));
    defparam \config_register_latched_dec_inst1.STATSR_29_LC_18_28_7 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_29_LC_18_28_7 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_29_LC_18_28_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_29_LC_18_28_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6240),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6184),
            .ce(N__5952),
            .sr(N__5866));
    defparam \config_register_latched_dec_inst1.STATSR_60_LC_18_30_0 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_60_LC_18_30_0 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_60_LC_18_30_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_60_LC_18_30_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6216),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6186),
            .ce(N__5946),
            .sr(N__5868));
    defparam \config_register_latched_dec_inst1.STATSR_55_LC_18_30_1 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_55_LC_18_30_1 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_55_LC_18_30_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_55_LC_18_30_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6222),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6186),
            .ce(N__5946),
            .sr(N__5868));
    defparam \config_register_latched_dec_inst1.STATSR_59_LC_18_30_2 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_59_LC_18_30_2 .SEQ_MODE=4'b1011;
    defparam \config_register_latched_dec_inst1.STATSR_59_LC_18_30_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_59_LC_18_30_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6204),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6186),
            .ce(N__5946),
            .sr(N__5868));
    defparam \config_register_latched_dec_inst1.STATSR_57_LC_18_30_3 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_57_LC_18_30_3 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_57_LC_18_30_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_57_LC_18_30_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6192),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6186),
            .ce(N__5946),
            .sr(N__5868));
    defparam \config_register_latched_dec_inst1.STATSR_58_LC_18_30_4 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_58_LC_18_30_4 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_58_LC_18_30_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_58_LC_18_30_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6210),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6186),
            .ce(N__5946),
            .sr(N__5868));
    defparam \config_register_latched_dec_inst1.STATSR_56_LC_18_30_6 .C_ON=1'b0;
    defparam \config_register_latched_dec_inst1.STATSR_56_LC_18_30_6 .SEQ_MODE=4'b1010;
    defparam \config_register_latched_dec_inst1.STATSR_56_LC_18_30_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \config_register_latched_dec_inst1.STATSR_56_LC_18_30_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6198),
            .lcout(\config_register_latched_dec_inst1.STATSRZ0Z_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6186),
            .ce(N__5946),
            .sr(N__5868));
endmodule // top
