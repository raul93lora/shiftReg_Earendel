// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 13 2025 09:41:53

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    signal_out,
    CLK,
    SELSTAT,
    SELDYN,
    RST_N);

    output signal_out;
    input CLK;
    input SELSTAT;
    input SELDYN;
    input RST_N;

    wire N__2336;
    wire N__2335;
    wire N__2334;
    wire N__2325;
    wire N__2324;
    wire N__2323;
    wire N__2316;
    wire N__2315;
    wire N__2314;
    wire N__2307;
    wire N__2306;
    wire N__2305;
    wire N__2298;
    wire N__2297;
    wire N__2296;
    wire N__2279;
    wire N__2276;
    wire N__2273;
    wire N__2270;
    wire N__2267;
    wire N__2264;
    wire N__2261;
    wire N__2258;
    wire N__2255;
    wire N__2252;
    wire N__2249;
    wire N__2246;
    wire N__2243;
    wire N__2240;
    wire N__2237;
    wire N__2234;
    wire N__2231;
    wire N__2228;
    wire N__2225;
    wire N__2222;
    wire N__2219;
    wire N__2216;
    wire N__2213;
    wire N__2210;
    wire N__2207;
    wire N__2206;
    wire N__2205;
    wire N__2204;
    wire N__2203;
    wire N__2202;
    wire N__2201;
    wire N__2200;
    wire N__2199;
    wire N__2198;
    wire N__2197;
    wire N__2196;
    wire N__2195;
    wire N__2194;
    wire N__2193;
    wire N__2192;
    wire N__2191;
    wire N__2156;
    wire N__2153;
    wire N__2150;
    wire N__2149;
    wire N__2148;
    wire N__2147;
    wire N__2146;
    wire N__2145;
    wire N__2144;
    wire N__2143;
    wire N__2142;
    wire N__2141;
    wire N__2140;
    wire N__2139;
    wire N__2138;
    wire N__2137;
    wire N__2108;
    wire N__2105;
    wire N__2102;
    wire N__2101;
    wire N__2100;
    wire N__2099;
    wire N__2098;
    wire N__2097;
    wire N__2096;
    wire N__2095;
    wire N__2094;
    wire N__2093;
    wire N__2092;
    wire N__2091;
    wire N__2090;
    wire N__2089;
    wire N__2088;
    wire N__2087;
    wire N__2086;
    wire N__2051;
    wire N__2048;
    wire N__2045;
    wire N__2042;
    wire N__2039;
    wire N__2036;
    wire N__2033;
    wire N__2030;
    wire N__2027;
    wire N__2024;
    wire N__2021;
    wire N__2018;
    wire N__2015;
    wire N__2012;
    wire N__2009;
    wire N__2006;
    wire N__2003;
    wire N__2000;
    wire N__1997;
    wire N__1994;
    wire N__1991;
    wire N__1988;
    wire N__1985;
    wire N__1982;
    wire N__1979;
    wire N__1976;
    wire N__1973;
    wire N__1970;
    wire N__1967;
    wire N__1964;
    wire N__1961;
    wire N__1958;
    wire N__1955;
    wire N__1952;
    wire N__1949;
    wire N__1946;
    wire N__1943;
    wire N__1940;
    wire N__1937;
    wire N__1934;
    wire N__1931;
    wire N__1928;
    wire N__1925;
    wire N__1922;
    wire N__1919;
    wire N__1916;
    wire N__1913;
    wire N__1910;
    wire N__1907;
    wire N__1904;
    wire N__1901;
    wire N__1898;
    wire N__1895;
    wire N__1892;
    wire N__1889;
    wire N__1886;
    wire N__1883;
    wire N__1880;
    wire N__1877;
    wire N__1874;
    wire N__1871;
    wire N__1868;
    wire N__1865;
    wire N__1862;
    wire N__1859;
    wire N__1856;
    wire N__1853;
    wire N__1850;
    wire N__1847;
    wire N__1844;
    wire N__1841;
    wire N__1838;
    wire N__1835;
    wire N__1832;
    wire N__1829;
    wire N__1826;
    wire N__1823;
    wire N__1820;
    wire N__1817;
    wire N__1814;
    wire N__1811;
    wire N__1808;
    wire N__1805;
    wire N__1802;
    wire N__1799;
    wire N__1796;
    wire N__1793;
    wire N__1790;
    wire N__1787;
    wire N__1784;
    wire N__1781;
    wire N__1778;
    wire N__1775;
    wire N__1772;
    wire N__1769;
    wire N__1766;
    wire N__1763;
    wire N__1760;
    wire N__1757;
    wire N__1754;
    wire N__1751;
    wire N__1748;
    wire N__1745;
    wire N__1742;
    wire N__1739;
    wire N__1736;
    wire N__1733;
    wire N__1730;
    wire N__1727;
    wire N__1724;
    wire N__1721;
    wire N__1718;
    wire N__1715;
    wire N__1712;
    wire N__1709;
    wire N__1706;
    wire N__1703;
    wire N__1700;
    wire N__1697;
    wire N__1694;
    wire N__1691;
    wire N__1688;
    wire N__1685;
    wire N__1682;
    wire N__1679;
    wire N__1676;
    wire N__1673;
    wire N__1670;
    wire N__1667;
    wire N__1664;
    wire N__1661;
    wire N__1658;
    wire N__1655;
    wire N__1652;
    wire N__1649;
    wire N__1646;
    wire N__1643;
    wire N__1640;
    wire N__1637;
    wire N__1634;
    wire N__1631;
    wire N__1628;
    wire N__1625;
    wire N__1622;
    wire N__1619;
    wire N__1616;
    wire N__1613;
    wire N__1610;
    wire N__1607;
    wire N__1604;
    wire N__1601;
    wire N__1598;
    wire N__1595;
    wire N__1592;
    wire N__1589;
    wire N__1586;
    wire N__1583;
    wire N__1580;
    wire N__1577;
    wire N__1574;
    wire N__1571;
    wire N__1570;
    wire N__1567;
    wire N__1564;
    wire N__1559;
    wire N__1556;
    wire N__1555;
    wire N__1552;
    wire N__1549;
    wire N__1544;
    wire N__1543;
    wire N__1540;
    wire N__1537;
    wire N__1536;
    wire N__1531;
    wire N__1528;
    wire N__1523;
    wire N__1520;
    wire N__1517;
    wire N__1514;
    wire N__1511;
    wire N__1508;
    wire N__1505;
    wire N__1502;
    wire N__1499;
    wire N__1496;
    wire N__1493;
    wire N__1490;
    wire N__1487;
    wire N__1484;
    wire N__1481;
    wire N__1478;
    wire N__1475;
    wire N__1472;
    wire N__1469;
    wire N__1466;
    wire N__1463;
    wire N__1460;
    wire N__1457;
    wire N__1454;
    wire N__1451;
    wire N__1448;
    wire N__1445;
    wire N__1442;
    wire N__1439;
    wire N__1436;
    wire N__1433;
    wire N__1430;
    wire N__1427;
    wire N__1424;
    wire N__1421;
    wire N__1418;
    wire N__1415;
    wire N__1412;
    wire N__1409;
    wire N__1406;
    wire N__1403;
    wire N__1400;
    wire N__1397;
    wire N__1394;
    wire N__1391;
    wire N__1388;
    wire N__1385;
    wire N__1382;
    wire N__1379;
    wire N__1376;
    wire N__1373;
    wire N__1370;
    wire VCCG0;
    wire RST_N_c;
    wire RST_N_c_i;
    wire generated_signal;
    wire signal_out_c;
    wire \generator_inst1.REGDYNZ0Z_8 ;
    wire \generator_inst1.REGDYNZ0Z_12 ;
    wire \generator_inst1.REGDYNZ0Z_13 ;
    wire \generator_inst1.REGDYNZ0Z_14 ;
    wire \generator_inst1.REGDYNZ0Z_15 ;
    wire \generator_inst1.REGDYNZ0Z_11 ;
    wire \generator_inst1.REGDYNZ0Z_9 ;
    wire \generator_inst1.REGDYNZ0Z_10 ;
    wire \generator_inst1.REGDYNZ0Z_1 ;
    wire \generator_inst1.REGDYNZ0Z_2 ;
    wire \generator_inst1.REGDYNZ0Z_6 ;
    wire \generator_inst1.REGDYNZ0Z_7 ;
    wire \generator_inst1.REGDYNZ0Z_5 ;
    wire \generator_inst1.REGDYNZ0Z_3 ;
    wire \generator_inst1.REGDYNZ0Z_4 ;
    wire \generator_inst1.REGDYNZ0Z_0 ;
    wire \generator_inst1.REGSTATZ0Z_24 ;
    wire \generator_inst1.REGSTATZ0Z_25 ;
    wire \generator_inst1.REGSTATZ0Z_22 ;
    wire \generator_inst1.REGSTATZ0Z_23 ;
    wire \generator_inst1.REGSTATZ0Z_21 ;
    wire SELSTAT_c;
    wire SELDYN_c;
    wire \generator_inst1.REGDYNZ0Z7 ;
    wire \generator_inst1.REGSTATZ0Z_83 ;
    wire \generator_inst1.REGSTATZ0Z_84 ;
    wire \generator_inst1.REGSTATZ0Z_87 ;
    wire \generator_inst1.REGSTATZ0Z_85 ;
    wire \generator_inst1.REGSTATZ0Z_86 ;
    wire \generator_inst1.REGSTATZ0Z_81 ;
    wire \generator_inst1.REGSTATZ0Z_82 ;
    wire \generator_inst1.REGSTATZ0Z_77 ;
    wire \generator_inst1.REGSTATZ0Z_78 ;
    wire \generator_inst1.REGSTATZ0Z_79 ;
    wire \generator_inst1.REGSTATZ0Z_80 ;
    wire \generator_inst1.REGSTATZ0Z_76 ;
    wire \generator_inst1.REGSTATZ0Z_73 ;
    wire \generator_inst1.REGSTATZ0Z_74 ;
    wire \generator_inst1.REGSTATZ0Z_75 ;
    wire \generator_inst1.REGSTATZ0Z_14 ;
    wire \generator_inst1.REGSTATZ0Z_17 ;
    wire \generator_inst1.REGSTATZ0Z_15 ;
    wire \generator_inst1.REGSTATZ0Z_16 ;
    wire \generator_inst1.REGSTATZ0Z_47 ;
    wire \generator_inst1.REGSTATZ0Z_48 ;
    wire \generator_inst1.REGSTATZ0Z_18 ;
    wire \generator_inst1.REGSTATZ0Z_19 ;
    wire \generator_inst1.REGSTATZ0Z_20 ;
    wire \generator_inst1.REGSTATZ0Z_28 ;
    wire \generator_inst1.REGSTATZ0Z_29 ;
    wire \generator_inst1.REGSTATZ0Z_30 ;
    wire \generator_inst1.REGSTATZ0Z_31 ;
    wire \generator_inst1.REGSTATZ0Z_32 ;
    wire \generator_inst1.REGSTATZ0Z_26 ;
    wire \generator_inst1.REGSTATZ0Z_27 ;
    wire \generator_inst1.REGSTATZ0Z_11 ;
    wire \generator_inst1.REGSTATZ0Z_6 ;
    wire \generator_inst1.REGSTATZ0Z_10 ;
    wire \generator_inst1.REGSTATZ0Z_7 ;
    wire \generator_inst1.REGSTATZ0Z_8 ;
    wire \generator_inst1.REGSTATZ0Z_9 ;
    wire \generator_inst1.REGSTATZ0Z_62 ;
    wire \generator_inst1.REGSTATZ0Z_63 ;
    wire \generator_inst1.REGSTATZ0Z_72 ;
    wire \generator_inst1.REGSTATZ0Z_60 ;
    wire \generator_inst1.REGSTATZ0Z_61 ;
    wire \generator_inst1.REGSTATZ0Z_12 ;
    wire \generator_inst1.REGSTATZ0Z_13 ;
    wire \generator_inst1.REGSTATZ0Z_64 ;
    wire \generator_inst1.REGSTATZ0Z_49 ;
    wire \generator_inst1.REGSTATZ0Z_50 ;
    wire \generator_inst1.REGSTATZ0Z_51 ;
    wire \generator_inst1.REGSTATZ0Z_54 ;
    wire \generator_inst1.REGSTATZ0Z_52 ;
    wire \generator_inst1.REGSTATZ0Z_53 ;
    wire \generator_inst1.REGSTATZ0Z_43 ;
    wire \generator_inst1.REGSTATZ0Z_44 ;
    wire \generator_inst1.REGSTATZ0Z_45 ;
    wire \generator_inst1.REGSTATZ0Z_46 ;
    wire \generator_inst1.REGSTATZ0Z_33 ;
    wire GNDG0;
    wire \generator_inst1.REGSTATZ0Z_2 ;
    wire \generator_inst1.REGSTATZ0Z_5 ;
    wire \generator_inst1.REGSTATZ0Z_0 ;
    wire \generator_inst1.REGSTATZ0Z_1 ;
    wire \generator_inst1.REGSTATZ0Z_3 ;
    wire \generator_inst1.REGSTATZ0Z_4 ;
    wire \generator_inst1.REGSTATZ0Z_65 ;
    wire \generator_inst1.REGSTATZ0Z_66 ;
    wire \generator_inst1.REGSTATZ0Z_71 ;
    wire \generator_inst1.REGSTATZ0Z_69 ;
    wire \generator_inst1.REGSTATZ0Z_70 ;
    wire \generator_inst1.REGSTATZ0Z_67 ;
    wire \generator_inst1.REGSTATZ0Z_68 ;
    wire \generator_inst1.REGSTATZ0Z_55 ;
    wire \generator_inst1.REGSTATZ0Z_56 ;
    wire \generator_inst1.REGSTATZ0Z_57 ;
    wire \generator_inst1.REGSTATZ0Z_58 ;
    wire \generator_inst1.REGSTATZ0Z_59 ;
    wire \generator_inst1.REGSTATZ0Z_36 ;
    wire \generator_inst1.REGSTATZ0Z_37 ;
    wire \generator_inst1.REGSTATZ0Z_38 ;
    wire \generator_inst1.REGSTATZ0Z_42 ;
    wire \generator_inst1.REGSTATZ0Z_39 ;
    wire \generator_inst1.REGSTATZ0Z_40 ;
    wire \generator_inst1.REGSTATZ0Z_41 ;
    wire \generator_inst1.REGSTATZ0Z_34 ;
    wire \generator_inst1.REGSTATZ0Z_35 ;
    wire _gnd_net_;
    wire CLK_c_g;
    wire \generator_inst1.REGDYN7_g ;
    wire RST_N_c_i_g;

    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__2334),
            .GLOBALBUFFEROUTPUT(CLK_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__2336),
            .DIN(N__2335),
            .DOUT(N__2334),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__2336),
            .PADOUT(N__2335),
            .PADIN(N__2334),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RST_N_ibuf_iopad (
            .OE(N__2325),
            .DIN(N__2324),
            .DOUT(N__2323),
            .PACKAGEPIN(RST_N));
    defparam RST_N_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RST_N_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RST_N_ibuf_preio (
            .PADOEN(N__2325),
            .PADOUT(N__2324),
            .PADIN(N__2323),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RST_N_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SELDYN_ibuf_iopad (
            .OE(N__2316),
            .DIN(N__2315),
            .DOUT(N__2314),
            .PACKAGEPIN(SELDYN));
    defparam SELDYN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SELDYN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SELDYN_ibuf_preio (
            .PADOEN(N__2316),
            .PADOUT(N__2315),
            .PADIN(N__2314),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SELDYN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD signal_out_obuf_iopad (
            .OE(N__2307),
            .DIN(N__2306),
            .DOUT(N__2305),
            .PACKAGEPIN(signal_out));
    defparam signal_out_obuf_preio.NEG_TRIGGER=1'b0;
    defparam signal_out_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO signal_out_obuf_preio (
            .PADOEN(N__2307),
            .PADOUT(N__2306),
            .PADIN(N__2305),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1418),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SELSTAT_ibuf_iopad (
            .OE(N__2298),
            .DIN(N__2297),
            .DOUT(N__2296),
            .PACKAGEPIN(SELSTAT));
    defparam SELSTAT_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SELSTAT_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SELSTAT_ibuf_preio (
            .PADOEN(N__2298),
            .PADOUT(N__2297),
            .PADIN(N__2296),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SELSTAT_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__421 (
            .O(N__2279),
            .I(N__2276));
    LocalMux I__420 (
            .O(N__2276),
            .I(\generator_inst1.REGSTATZ0Z_57 ));
    InMux I__419 (
            .O(N__2273),
            .I(N__2270));
    LocalMux I__418 (
            .O(N__2270),
            .I(\generator_inst1.REGSTATZ0Z_58 ));
    InMux I__417 (
            .O(N__2267),
            .I(N__2264));
    LocalMux I__416 (
            .O(N__2264),
            .I(\generator_inst1.REGSTATZ0Z_59 ));
    InMux I__415 (
            .O(N__2261),
            .I(N__2258));
    LocalMux I__414 (
            .O(N__2258),
            .I(\generator_inst1.REGSTATZ0Z_36 ));
    InMux I__413 (
            .O(N__2255),
            .I(N__2252));
    LocalMux I__412 (
            .O(N__2252),
            .I(\generator_inst1.REGSTATZ0Z_37 ));
    InMux I__411 (
            .O(N__2249),
            .I(N__2246));
    LocalMux I__410 (
            .O(N__2246),
            .I(\generator_inst1.REGSTATZ0Z_38 ));
    InMux I__409 (
            .O(N__2243),
            .I(N__2240));
    LocalMux I__408 (
            .O(N__2240),
            .I(\generator_inst1.REGSTATZ0Z_42 ));
    InMux I__407 (
            .O(N__2237),
            .I(N__2234));
    LocalMux I__406 (
            .O(N__2234),
            .I(\generator_inst1.REGSTATZ0Z_39 ));
    InMux I__405 (
            .O(N__2231),
            .I(N__2228));
    LocalMux I__404 (
            .O(N__2228),
            .I(\generator_inst1.REGSTATZ0Z_40 ));
    InMux I__403 (
            .O(N__2225),
            .I(N__2222));
    LocalMux I__402 (
            .O(N__2222),
            .I(\generator_inst1.REGSTATZ0Z_41 ));
    InMux I__401 (
            .O(N__2219),
            .I(N__2216));
    LocalMux I__400 (
            .O(N__2216),
            .I(\generator_inst1.REGSTATZ0Z_34 ));
    InMux I__399 (
            .O(N__2213),
            .I(N__2210));
    LocalMux I__398 (
            .O(N__2210),
            .I(\generator_inst1.REGSTATZ0Z_35 ));
    ClkMux I__397 (
            .O(N__2207),
            .I(N__2156));
    ClkMux I__396 (
            .O(N__2206),
            .I(N__2156));
    ClkMux I__395 (
            .O(N__2205),
            .I(N__2156));
    ClkMux I__394 (
            .O(N__2204),
            .I(N__2156));
    ClkMux I__393 (
            .O(N__2203),
            .I(N__2156));
    ClkMux I__392 (
            .O(N__2202),
            .I(N__2156));
    ClkMux I__391 (
            .O(N__2201),
            .I(N__2156));
    ClkMux I__390 (
            .O(N__2200),
            .I(N__2156));
    ClkMux I__389 (
            .O(N__2199),
            .I(N__2156));
    ClkMux I__388 (
            .O(N__2198),
            .I(N__2156));
    ClkMux I__387 (
            .O(N__2197),
            .I(N__2156));
    ClkMux I__386 (
            .O(N__2196),
            .I(N__2156));
    ClkMux I__385 (
            .O(N__2195),
            .I(N__2156));
    ClkMux I__384 (
            .O(N__2194),
            .I(N__2156));
    ClkMux I__383 (
            .O(N__2193),
            .I(N__2156));
    ClkMux I__382 (
            .O(N__2192),
            .I(N__2156));
    ClkMux I__381 (
            .O(N__2191),
            .I(N__2156));
    GlobalMux I__380 (
            .O(N__2156),
            .I(N__2153));
    gio2CtrlBuf I__379 (
            .O(N__2153),
            .I(CLK_c_g));
    CEMux I__378 (
            .O(N__2150),
            .I(N__2108));
    CEMux I__377 (
            .O(N__2149),
            .I(N__2108));
    CEMux I__376 (
            .O(N__2148),
            .I(N__2108));
    CEMux I__375 (
            .O(N__2147),
            .I(N__2108));
    CEMux I__374 (
            .O(N__2146),
            .I(N__2108));
    CEMux I__373 (
            .O(N__2145),
            .I(N__2108));
    CEMux I__372 (
            .O(N__2144),
            .I(N__2108));
    CEMux I__371 (
            .O(N__2143),
            .I(N__2108));
    CEMux I__370 (
            .O(N__2142),
            .I(N__2108));
    CEMux I__369 (
            .O(N__2141),
            .I(N__2108));
    CEMux I__368 (
            .O(N__2140),
            .I(N__2108));
    CEMux I__367 (
            .O(N__2139),
            .I(N__2108));
    CEMux I__366 (
            .O(N__2138),
            .I(N__2108));
    CEMux I__365 (
            .O(N__2137),
            .I(N__2108));
    GlobalMux I__364 (
            .O(N__2108),
            .I(N__2105));
    gio2CtrlBuf I__363 (
            .O(N__2105),
            .I(\generator_inst1.REGDYN7_g ));
    SRMux I__362 (
            .O(N__2102),
            .I(N__2051));
    SRMux I__361 (
            .O(N__2101),
            .I(N__2051));
    SRMux I__360 (
            .O(N__2100),
            .I(N__2051));
    SRMux I__359 (
            .O(N__2099),
            .I(N__2051));
    SRMux I__358 (
            .O(N__2098),
            .I(N__2051));
    SRMux I__357 (
            .O(N__2097),
            .I(N__2051));
    SRMux I__356 (
            .O(N__2096),
            .I(N__2051));
    SRMux I__355 (
            .O(N__2095),
            .I(N__2051));
    SRMux I__354 (
            .O(N__2094),
            .I(N__2051));
    SRMux I__353 (
            .O(N__2093),
            .I(N__2051));
    SRMux I__352 (
            .O(N__2092),
            .I(N__2051));
    SRMux I__351 (
            .O(N__2091),
            .I(N__2051));
    SRMux I__350 (
            .O(N__2090),
            .I(N__2051));
    SRMux I__349 (
            .O(N__2089),
            .I(N__2051));
    SRMux I__348 (
            .O(N__2088),
            .I(N__2051));
    SRMux I__347 (
            .O(N__2087),
            .I(N__2051));
    SRMux I__346 (
            .O(N__2086),
            .I(N__2051));
    GlobalMux I__345 (
            .O(N__2051),
            .I(N__2048));
    gio2CtrlBuf I__344 (
            .O(N__2048),
            .I(RST_N_c_i_g));
    InMux I__343 (
            .O(N__2045),
            .I(N__2042));
    LocalMux I__342 (
            .O(N__2042),
            .I(\generator_inst1.REGSTATZ0Z_66 ));
    InMux I__341 (
            .O(N__2039),
            .I(N__2036));
    LocalMux I__340 (
            .O(N__2036),
            .I(\generator_inst1.REGSTATZ0Z_71 ));
    InMux I__339 (
            .O(N__2033),
            .I(N__2030));
    LocalMux I__338 (
            .O(N__2030),
            .I(\generator_inst1.REGSTATZ0Z_69 ));
    InMux I__337 (
            .O(N__2027),
            .I(N__2024));
    LocalMux I__336 (
            .O(N__2024),
            .I(\generator_inst1.REGSTATZ0Z_70 ));
    InMux I__335 (
            .O(N__2021),
            .I(N__2018));
    LocalMux I__334 (
            .O(N__2018),
            .I(\generator_inst1.REGSTATZ0Z_67 ));
    InMux I__333 (
            .O(N__2015),
            .I(N__2012));
    LocalMux I__332 (
            .O(N__2012),
            .I(\generator_inst1.REGSTATZ0Z_68 ));
    InMux I__331 (
            .O(N__2009),
            .I(N__2006));
    LocalMux I__330 (
            .O(N__2006),
            .I(\generator_inst1.REGSTATZ0Z_55 ));
    InMux I__329 (
            .O(N__2003),
            .I(N__2000));
    LocalMux I__328 (
            .O(N__2000),
            .I(\generator_inst1.REGSTATZ0Z_56 ));
    InMux I__327 (
            .O(N__1997),
            .I(N__1994));
    LocalMux I__326 (
            .O(N__1994),
            .I(\generator_inst1.REGSTATZ0Z_45 ));
    InMux I__325 (
            .O(N__1991),
            .I(N__1988));
    LocalMux I__324 (
            .O(N__1988),
            .I(\generator_inst1.REGSTATZ0Z_46 ));
    InMux I__323 (
            .O(N__1985),
            .I(N__1982));
    LocalMux I__322 (
            .O(N__1982),
            .I(\generator_inst1.REGSTATZ0Z_33 ));
    InMux I__321 (
            .O(N__1979),
            .I(N__1976));
    LocalMux I__320 (
            .O(N__1976),
            .I(\generator_inst1.REGSTATZ0Z_2 ));
    InMux I__319 (
            .O(N__1973),
            .I(N__1970));
    LocalMux I__318 (
            .O(N__1970),
            .I(\generator_inst1.REGSTATZ0Z_5 ));
    InMux I__317 (
            .O(N__1967),
            .I(N__1964));
    LocalMux I__316 (
            .O(N__1964),
            .I(\generator_inst1.REGSTATZ0Z_0 ));
    InMux I__315 (
            .O(N__1961),
            .I(N__1958));
    LocalMux I__314 (
            .O(N__1958),
            .I(\generator_inst1.REGSTATZ0Z_1 ));
    InMux I__313 (
            .O(N__1955),
            .I(N__1952));
    LocalMux I__312 (
            .O(N__1952),
            .I(\generator_inst1.REGSTATZ0Z_3 ));
    InMux I__311 (
            .O(N__1949),
            .I(N__1946));
    LocalMux I__310 (
            .O(N__1946),
            .I(\generator_inst1.REGSTATZ0Z_4 ));
    InMux I__309 (
            .O(N__1943),
            .I(N__1940));
    LocalMux I__308 (
            .O(N__1940),
            .I(\generator_inst1.REGSTATZ0Z_65 ));
    InMux I__307 (
            .O(N__1937),
            .I(N__1934));
    LocalMux I__306 (
            .O(N__1934),
            .I(\generator_inst1.REGSTATZ0Z_49 ));
    InMux I__305 (
            .O(N__1931),
            .I(N__1928));
    LocalMux I__304 (
            .O(N__1928),
            .I(\generator_inst1.REGSTATZ0Z_50 ));
    InMux I__303 (
            .O(N__1925),
            .I(N__1922));
    LocalMux I__302 (
            .O(N__1922),
            .I(\generator_inst1.REGSTATZ0Z_51 ));
    InMux I__301 (
            .O(N__1919),
            .I(N__1916));
    LocalMux I__300 (
            .O(N__1916),
            .I(\generator_inst1.REGSTATZ0Z_54 ));
    InMux I__299 (
            .O(N__1913),
            .I(N__1910));
    LocalMux I__298 (
            .O(N__1910),
            .I(\generator_inst1.REGSTATZ0Z_52 ));
    InMux I__297 (
            .O(N__1907),
            .I(N__1904));
    LocalMux I__296 (
            .O(N__1904),
            .I(\generator_inst1.REGSTATZ0Z_53 ));
    InMux I__295 (
            .O(N__1901),
            .I(N__1898));
    LocalMux I__294 (
            .O(N__1898),
            .I(\generator_inst1.REGSTATZ0Z_43 ));
    InMux I__293 (
            .O(N__1895),
            .I(N__1892));
    LocalMux I__292 (
            .O(N__1892),
            .I(\generator_inst1.REGSTATZ0Z_44 ));
    InMux I__291 (
            .O(N__1889),
            .I(N__1886));
    LocalMux I__290 (
            .O(N__1886),
            .I(\generator_inst1.REGSTATZ0Z_8 ));
    InMux I__289 (
            .O(N__1883),
            .I(N__1880));
    LocalMux I__288 (
            .O(N__1880),
            .I(\generator_inst1.REGSTATZ0Z_9 ));
    InMux I__287 (
            .O(N__1877),
            .I(N__1874));
    LocalMux I__286 (
            .O(N__1874),
            .I(\generator_inst1.REGSTATZ0Z_62 ));
    InMux I__285 (
            .O(N__1871),
            .I(N__1868));
    LocalMux I__284 (
            .O(N__1868),
            .I(\generator_inst1.REGSTATZ0Z_63 ));
    InMux I__283 (
            .O(N__1865),
            .I(N__1862));
    LocalMux I__282 (
            .O(N__1862),
            .I(\generator_inst1.REGSTATZ0Z_72 ));
    InMux I__281 (
            .O(N__1859),
            .I(N__1856));
    LocalMux I__280 (
            .O(N__1856),
            .I(\generator_inst1.REGSTATZ0Z_60 ));
    InMux I__279 (
            .O(N__1853),
            .I(N__1850));
    LocalMux I__278 (
            .O(N__1850),
            .I(\generator_inst1.REGSTATZ0Z_61 ));
    CascadeMux I__277 (
            .O(N__1847),
            .I(N__1844));
    InMux I__276 (
            .O(N__1844),
            .I(N__1841));
    LocalMux I__275 (
            .O(N__1841),
            .I(\generator_inst1.REGSTATZ0Z_12 ));
    InMux I__274 (
            .O(N__1838),
            .I(N__1835));
    LocalMux I__273 (
            .O(N__1835),
            .I(\generator_inst1.REGSTATZ0Z_13 ));
    InMux I__272 (
            .O(N__1832),
            .I(N__1829));
    LocalMux I__271 (
            .O(N__1829),
            .I(\generator_inst1.REGSTATZ0Z_64 ));
    InMux I__270 (
            .O(N__1826),
            .I(N__1823));
    LocalMux I__269 (
            .O(N__1823),
            .I(\generator_inst1.REGSTATZ0Z_30 ));
    InMux I__268 (
            .O(N__1820),
            .I(N__1817));
    LocalMux I__267 (
            .O(N__1817),
            .I(\generator_inst1.REGSTATZ0Z_31 ));
    InMux I__266 (
            .O(N__1814),
            .I(N__1811));
    LocalMux I__265 (
            .O(N__1811),
            .I(\generator_inst1.REGSTATZ0Z_32 ));
    InMux I__264 (
            .O(N__1808),
            .I(N__1805));
    LocalMux I__263 (
            .O(N__1805),
            .I(\generator_inst1.REGSTATZ0Z_26 ));
    InMux I__262 (
            .O(N__1802),
            .I(N__1799));
    LocalMux I__261 (
            .O(N__1799),
            .I(\generator_inst1.REGSTATZ0Z_27 ));
    InMux I__260 (
            .O(N__1796),
            .I(N__1793));
    LocalMux I__259 (
            .O(N__1793),
            .I(\generator_inst1.REGSTATZ0Z_11 ));
    InMux I__258 (
            .O(N__1790),
            .I(N__1787));
    LocalMux I__257 (
            .O(N__1787),
            .I(\generator_inst1.REGSTATZ0Z_6 ));
    InMux I__256 (
            .O(N__1784),
            .I(N__1781));
    LocalMux I__255 (
            .O(N__1781),
            .I(\generator_inst1.REGSTATZ0Z_10 ));
    InMux I__254 (
            .O(N__1778),
            .I(N__1775));
    LocalMux I__253 (
            .O(N__1775),
            .I(\generator_inst1.REGSTATZ0Z_7 ));
    CascadeMux I__252 (
            .O(N__1772),
            .I(N__1769));
    InMux I__251 (
            .O(N__1769),
            .I(N__1766));
    LocalMux I__250 (
            .O(N__1766),
            .I(\generator_inst1.REGSTATZ0Z_15 ));
    InMux I__249 (
            .O(N__1763),
            .I(N__1760));
    LocalMux I__248 (
            .O(N__1760),
            .I(\generator_inst1.REGSTATZ0Z_16 ));
    InMux I__247 (
            .O(N__1757),
            .I(N__1754));
    LocalMux I__246 (
            .O(N__1754),
            .I(\generator_inst1.REGSTATZ0Z_47 ));
    InMux I__245 (
            .O(N__1751),
            .I(N__1748));
    LocalMux I__244 (
            .O(N__1748),
            .I(\generator_inst1.REGSTATZ0Z_48 ));
    InMux I__243 (
            .O(N__1745),
            .I(N__1742));
    LocalMux I__242 (
            .O(N__1742),
            .I(\generator_inst1.REGSTATZ0Z_18 ));
    InMux I__241 (
            .O(N__1739),
            .I(N__1736));
    LocalMux I__240 (
            .O(N__1736),
            .I(\generator_inst1.REGSTATZ0Z_19 ));
    InMux I__239 (
            .O(N__1733),
            .I(N__1730));
    LocalMux I__238 (
            .O(N__1730),
            .I(\generator_inst1.REGSTATZ0Z_20 ));
    InMux I__237 (
            .O(N__1727),
            .I(N__1724));
    LocalMux I__236 (
            .O(N__1724),
            .I(\generator_inst1.REGSTATZ0Z_28 ));
    InMux I__235 (
            .O(N__1721),
            .I(N__1718));
    LocalMux I__234 (
            .O(N__1718),
            .I(\generator_inst1.REGSTATZ0Z_29 ));
    InMux I__233 (
            .O(N__1715),
            .I(N__1712));
    LocalMux I__232 (
            .O(N__1712),
            .I(\generator_inst1.REGSTATZ0Z_79 ));
    InMux I__231 (
            .O(N__1709),
            .I(N__1706));
    LocalMux I__230 (
            .O(N__1706),
            .I(\generator_inst1.REGSTATZ0Z_80 ));
    InMux I__229 (
            .O(N__1703),
            .I(N__1700));
    LocalMux I__228 (
            .O(N__1700),
            .I(\generator_inst1.REGSTATZ0Z_76 ));
    InMux I__227 (
            .O(N__1697),
            .I(N__1694));
    LocalMux I__226 (
            .O(N__1694),
            .I(\generator_inst1.REGSTATZ0Z_73 ));
    InMux I__225 (
            .O(N__1691),
            .I(N__1688));
    LocalMux I__224 (
            .O(N__1688),
            .I(\generator_inst1.REGSTATZ0Z_74 ));
    InMux I__223 (
            .O(N__1685),
            .I(N__1682));
    LocalMux I__222 (
            .O(N__1682),
            .I(\generator_inst1.REGSTATZ0Z_75 ));
    InMux I__221 (
            .O(N__1679),
            .I(N__1676));
    LocalMux I__220 (
            .O(N__1676),
            .I(\generator_inst1.REGSTATZ0Z_14 ));
    InMux I__219 (
            .O(N__1673),
            .I(N__1670));
    LocalMux I__218 (
            .O(N__1670),
            .I(\generator_inst1.REGSTATZ0Z_17 ));
    InMux I__217 (
            .O(N__1667),
            .I(N__1664));
    LocalMux I__216 (
            .O(N__1664),
            .I(\generator_inst1.REGSTATZ0Z_83 ));
    InMux I__215 (
            .O(N__1661),
            .I(N__1658));
    LocalMux I__214 (
            .O(N__1658),
            .I(\generator_inst1.REGSTATZ0Z_84 ));
    InMux I__213 (
            .O(N__1655),
            .I(N__1652));
    LocalMux I__212 (
            .O(N__1652),
            .I(\generator_inst1.REGSTATZ0Z_87 ));
    InMux I__211 (
            .O(N__1649),
            .I(N__1646));
    LocalMux I__210 (
            .O(N__1646),
            .I(\generator_inst1.REGSTATZ0Z_85 ));
    InMux I__209 (
            .O(N__1643),
            .I(N__1640));
    LocalMux I__208 (
            .O(N__1640),
            .I(\generator_inst1.REGSTATZ0Z_86 ));
    InMux I__207 (
            .O(N__1637),
            .I(N__1634));
    LocalMux I__206 (
            .O(N__1634),
            .I(\generator_inst1.REGSTATZ0Z_81 ));
    InMux I__205 (
            .O(N__1631),
            .I(N__1628));
    LocalMux I__204 (
            .O(N__1628),
            .I(\generator_inst1.REGSTATZ0Z_82 ));
    InMux I__203 (
            .O(N__1625),
            .I(N__1622));
    LocalMux I__202 (
            .O(N__1622),
            .I(\generator_inst1.REGSTATZ0Z_77 ));
    InMux I__201 (
            .O(N__1619),
            .I(N__1616));
    LocalMux I__200 (
            .O(N__1616),
            .I(\generator_inst1.REGSTATZ0Z_78 ));
    InMux I__199 (
            .O(N__1613),
            .I(N__1610));
    LocalMux I__198 (
            .O(N__1610),
            .I(\generator_inst1.REGDYNZ0Z_0 ));
    InMux I__197 (
            .O(N__1607),
            .I(N__1604));
    LocalMux I__196 (
            .O(N__1604),
            .I(\generator_inst1.REGSTATZ0Z_24 ));
    InMux I__195 (
            .O(N__1601),
            .I(N__1598));
    LocalMux I__194 (
            .O(N__1598),
            .I(\generator_inst1.REGSTATZ0Z_25 ));
    InMux I__193 (
            .O(N__1595),
            .I(N__1592));
    LocalMux I__192 (
            .O(N__1592),
            .I(\generator_inst1.REGSTATZ0Z_22 ));
    InMux I__191 (
            .O(N__1589),
            .I(N__1586));
    LocalMux I__190 (
            .O(N__1586),
            .I(\generator_inst1.REGSTATZ0Z_23 ));
    InMux I__189 (
            .O(N__1583),
            .I(N__1580));
    LocalMux I__188 (
            .O(N__1580),
            .I(\generator_inst1.REGSTATZ0Z_21 ));
    InMux I__187 (
            .O(N__1577),
            .I(N__1574));
    LocalMux I__186 (
            .O(N__1574),
            .I(N__1571));
    IoSpan4Mux I__185 (
            .O(N__1571),
            .I(N__1567));
    InMux I__184 (
            .O(N__1570),
            .I(N__1564));
    Odrv4 I__183 (
            .O(N__1567),
            .I(SELSTAT_c));
    LocalMux I__182 (
            .O(N__1564),
            .I(SELSTAT_c));
    InMux I__181 (
            .O(N__1559),
            .I(N__1556));
    LocalMux I__180 (
            .O(N__1556),
            .I(N__1552));
    CEMux I__179 (
            .O(N__1555),
            .I(N__1549));
    Span4Mux_h I__178 (
            .O(N__1552),
            .I(N__1544));
    LocalMux I__177 (
            .O(N__1549),
            .I(N__1544));
    Span4Mux_v I__176 (
            .O(N__1544),
            .I(N__1540));
    CEMux I__175 (
            .O(N__1543),
            .I(N__1537));
    Span4Mux_v I__174 (
            .O(N__1540),
            .I(N__1531));
    LocalMux I__173 (
            .O(N__1537),
            .I(N__1531));
    InMux I__172 (
            .O(N__1536),
            .I(N__1528));
    Span4Mux_v I__171 (
            .O(N__1531),
            .I(N__1523));
    LocalMux I__170 (
            .O(N__1528),
            .I(N__1523));
    Span4Mux_v I__169 (
            .O(N__1523),
            .I(N__1520));
    Odrv4 I__168 (
            .O(N__1520),
            .I(SELDYN_c));
    IoInMux I__167 (
            .O(N__1517),
            .I(N__1514));
    LocalMux I__166 (
            .O(N__1514),
            .I(\generator_inst1.REGDYNZ0Z7 ));
    InMux I__165 (
            .O(N__1511),
            .I(N__1508));
    LocalMux I__164 (
            .O(N__1508),
            .I(\generator_inst1.REGDYNZ0Z_11 ));
    InMux I__163 (
            .O(N__1505),
            .I(N__1502));
    LocalMux I__162 (
            .O(N__1502),
            .I(\generator_inst1.REGDYNZ0Z_9 ));
    InMux I__161 (
            .O(N__1499),
            .I(N__1496));
    LocalMux I__160 (
            .O(N__1496),
            .I(\generator_inst1.REGDYNZ0Z_10 ));
    InMux I__159 (
            .O(N__1493),
            .I(N__1490));
    LocalMux I__158 (
            .O(N__1490),
            .I(\generator_inst1.REGDYNZ0Z_1 ));
    InMux I__157 (
            .O(N__1487),
            .I(N__1484));
    LocalMux I__156 (
            .O(N__1484),
            .I(\generator_inst1.REGDYNZ0Z_2 ));
    InMux I__155 (
            .O(N__1481),
            .I(N__1478));
    LocalMux I__154 (
            .O(N__1478),
            .I(\generator_inst1.REGDYNZ0Z_6 ));
    InMux I__153 (
            .O(N__1475),
            .I(N__1472));
    LocalMux I__152 (
            .O(N__1472),
            .I(\generator_inst1.REGDYNZ0Z_7 ));
    InMux I__151 (
            .O(N__1469),
            .I(N__1466));
    LocalMux I__150 (
            .O(N__1466),
            .I(\generator_inst1.REGDYNZ0Z_5 ));
    InMux I__149 (
            .O(N__1463),
            .I(N__1460));
    LocalMux I__148 (
            .O(N__1460),
            .I(\generator_inst1.REGDYNZ0Z_3 ));
    InMux I__147 (
            .O(N__1457),
            .I(N__1454));
    LocalMux I__146 (
            .O(N__1454),
            .I(\generator_inst1.REGDYNZ0Z_4 ));
    InMux I__145 (
            .O(N__1451),
            .I(N__1448));
    LocalMux I__144 (
            .O(N__1448),
            .I(N__1445));
    Span4Mux_v I__143 (
            .O(N__1445),
            .I(N__1442));
    Odrv4 I__142 (
            .O(N__1442),
            .I(RST_N_c));
    IoInMux I__141 (
            .O(N__1439),
            .I(N__1436));
    LocalMux I__140 (
            .O(N__1436),
            .I(N__1433));
    Span4Mux_s0_h I__139 (
            .O(N__1433),
            .I(N__1430));
    Span4Mux_v I__138 (
            .O(N__1430),
            .I(N__1427));
    Odrv4 I__137 (
            .O(N__1427),
            .I(RST_N_c_i));
    InMux I__136 (
            .O(N__1424),
            .I(N__1421));
    LocalMux I__135 (
            .O(N__1421),
            .I(generated_signal));
    IoInMux I__134 (
            .O(N__1418),
            .I(N__1415));
    LocalMux I__133 (
            .O(N__1415),
            .I(N__1412));
    IoSpan4Mux I__132 (
            .O(N__1412),
            .I(N__1409));
    IoSpan4Mux I__131 (
            .O(N__1409),
            .I(N__1406));
    IoSpan4Mux I__130 (
            .O(N__1406),
            .I(N__1403));
    Odrv4 I__129 (
            .O(N__1403),
            .I(signal_out_c));
    InMux I__128 (
            .O(N__1400),
            .I(N__1397));
    LocalMux I__127 (
            .O(N__1397),
            .I(\generator_inst1.REGDYNZ0Z_8 ));
    InMux I__126 (
            .O(N__1394),
            .I(N__1391));
    LocalMux I__125 (
            .O(N__1391),
            .I(\generator_inst1.REGDYNZ0Z_12 ));
    InMux I__124 (
            .O(N__1388),
            .I(N__1385));
    LocalMux I__123 (
            .O(N__1385),
            .I(\generator_inst1.REGDYNZ0Z_13 ));
    InMux I__122 (
            .O(N__1382),
            .I(N__1379));
    LocalMux I__121 (
            .O(N__1379),
            .I(\generator_inst1.REGDYNZ0Z_14 ));
    CascadeMux I__120 (
            .O(N__1376),
            .I(N__1373));
    InMux I__119 (
            .O(N__1373),
            .I(N__1370));
    LocalMux I__118 (
            .O(N__1370),
            .I(\generator_inst1.REGDYNZ0Z_15 ));
    GND GND (
            .Y(GNDG0));
    ICE_GB \generator_inst1.REGDYN7_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__1517),
            .GLOBALBUFFEROUTPUT(\generator_inst1.REGDYN7_g ));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB RST_N_ibuf_RNIBJGC_0 (
            .USERSIGNALTOGLOBALBUFFER(N__1439),
            .GLOBALBUFFEROUTPUT(RST_N_c_i_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam RST_N_ibuf_RNIBJGC_LC_1_10_0.C_ON=1'b0;
    defparam RST_N_ibuf_RNIBJGC_LC_1_10_0.SEQ_MODE=4'b0000;
    defparam RST_N_ibuf_RNIBJGC_LC_1_10_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 RST_N_ibuf_RNIBJGC_LC_1_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1451),
            .lcout(RST_N_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.signal_out_LC_1_12_0 .C_ON=1'b0;
    defparam \generator_inst1.signal_out_LC_1_12_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.signal_out_LC_1_12_0 .LUT_INIT=16'b0110010000100000;
    LogicCell40 \generator_inst1.signal_out_LC_1_12_0  (
            .in0(N__1577),
            .in1(N__1559),
            .in2(N__1376),
            .in3(N__1655),
            .lcout(generated_signal),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2200),
            .ce(),
            .sr(N__2095));
    defparam \receptor_inst1.signal_out_LC_1_12_1 .C_ON=1'b0;
    defparam \receptor_inst1.signal_out_LC_1_12_1 .SEQ_MODE=4'b1010;
    defparam \receptor_inst1.signal_out_LC_1_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \receptor_inst1.signal_out_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1424),
            .lcout(signal_out_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2200),
            .ce(),
            .sr(N__2095));
    defparam \generator_inst1.REGDYN_9_LC_1_13_0 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_9_LC_1_13_0 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_9_LC_1_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGDYN_9_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1400),
            .lcout(\generator_inst1.REGDYNZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2196),
            .ce(N__1555),
            .sr(N__2092));
    defparam \generator_inst1.REGDYN_8_LC_1_13_1 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_8_LC_1_13_1 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_8_LC_1_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGDYN_8_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1475),
            .lcout(\generator_inst1.REGDYNZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2196),
            .ce(N__1555),
            .sr(N__2092));
    defparam \generator_inst1.REGDYN_12_LC_1_13_2 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_12_LC_1_13_2 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGDYN_12_LC_1_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGDYN_12_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1511),
            .lcout(\generator_inst1.REGDYNZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2196),
            .ce(N__1555),
            .sr(N__2092));
    defparam \generator_inst1.REGDYN_13_LC_1_13_3 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_13_LC_1_13_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_13_LC_1_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGDYN_13_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1394),
            .lcout(\generator_inst1.REGDYNZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2196),
            .ce(N__1555),
            .sr(N__2092));
    defparam \generator_inst1.REGDYN_14_LC_1_13_4 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_14_LC_1_13_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGDYN_14_LC_1_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGDYN_14_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1388),
            .lcout(\generator_inst1.REGDYNZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2196),
            .ce(N__1555),
            .sr(N__2092));
    defparam \generator_inst1.REGDYN_15_LC_1_13_5 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_15_LC_1_13_5 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_15_LC_1_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGDYN_15_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1382),
            .lcout(\generator_inst1.REGDYNZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2196),
            .ce(N__1555),
            .sr(N__2092));
    defparam \generator_inst1.REGDYN_11_LC_1_13_6 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_11_LC_1_13_6 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_11_LC_1_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGDYN_11_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1499),
            .lcout(\generator_inst1.REGDYNZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2196),
            .ce(N__1555),
            .sr(N__2092));
    defparam \generator_inst1.REGDYN_10_LC_1_13_7 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_10_LC_1_13_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGDYN_10_LC_1_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGDYN_10_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1505),
            .lcout(\generator_inst1.REGDYNZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2196),
            .ce(N__1555),
            .sr(N__2092));
    defparam \generator_inst1.REGDYN_1_LC_1_14_0 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_1_LC_1_14_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGDYN_1_LC_1_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGDYN_1_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1613),
            .lcout(\generator_inst1.REGDYNZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2193),
            .ce(N__1543),
            .sr(N__2089));
    defparam \generator_inst1.REGDYN_2_LC_1_14_1 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_2_LC_1_14_1 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_2_LC_1_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGDYN_2_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1493),
            .lcout(\generator_inst1.REGDYNZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2193),
            .ce(N__1543),
            .sr(N__2089));
    defparam \generator_inst1.REGDYN_3_LC_1_14_2 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_3_LC_1_14_2 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_3_LC_1_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGDYN_3_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1487),
            .lcout(\generator_inst1.REGDYNZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2193),
            .ce(N__1543),
            .sr(N__2089));
    defparam \generator_inst1.REGDYN_6_LC_1_14_3 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_6_LC_1_14_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_6_LC_1_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGDYN_6_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1469),
            .lcout(\generator_inst1.REGDYNZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2193),
            .ce(N__1543),
            .sr(N__2089));
    defparam \generator_inst1.REGDYN_7_LC_1_14_4 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_7_LC_1_14_4 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_7_LC_1_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGDYN_7_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1481),
            .lcout(\generator_inst1.REGDYNZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2193),
            .ce(N__1543),
            .sr(N__2089));
    defparam \generator_inst1.REGDYN_5_LC_1_14_5 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_5_LC_1_14_5 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGDYN_5_LC_1_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGDYN_5_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1457),
            .lcout(\generator_inst1.REGDYNZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2193),
            .ce(N__1543),
            .sr(N__2089));
    defparam \generator_inst1.REGDYN_4_LC_1_14_6 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_4_LC_1_14_6 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGDYN_4_LC_1_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGDYN_4_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1463),
            .lcout(\generator_inst1.REGDYNZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2193),
            .ce(N__1543),
            .sr(N__2089));
    defparam \generator_inst1.REGDYN_0_LC_1_14_7 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN_0_LC_1_14_7 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGDYN_0_LC_1_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGDYN_0_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\generator_inst1.REGDYNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2193),
            .ce(N__1543),
            .sr(N__2089));
    defparam \generator_inst1.REGSTAT_24_LC_1_15_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_24_LC_1_15_0 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_24_LC_1_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_24_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1589),
            .lcout(\generator_inst1.REGSTATZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2191),
            .ce(N__2137),
            .sr(N__2087));
    defparam \generator_inst1.REGSTAT_26_LC_1_15_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_26_LC_1_15_2 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_26_LC_1_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_26_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1601),
            .lcout(\generator_inst1.REGSTATZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2191),
            .ce(N__2137),
            .sr(N__2087));
    defparam \generator_inst1.REGSTAT_25_LC_1_15_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_25_LC_1_15_3 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_25_LC_1_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_25_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1607),
            .lcout(\generator_inst1.REGSTATZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2191),
            .ce(N__2137),
            .sr(N__2087));
    defparam \generator_inst1.REGSTAT_22_LC_1_15_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_22_LC_1_15_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_22_LC_1_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_22_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1583),
            .lcout(\generator_inst1.REGSTATZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2191),
            .ce(N__2137),
            .sr(N__2087));
    defparam \generator_inst1.REGSTAT_23_LC_1_15_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_23_LC_1_15_5 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_23_LC_1_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_23_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1595),
            .lcout(\generator_inst1.REGSTATZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2191),
            .ce(N__2137),
            .sr(N__2087));
    defparam \generator_inst1.REGSTAT_21_LC_1_15_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_21_LC_1_15_7 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_21_LC_1_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_21_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1733),
            .lcout(\generator_inst1.REGSTATZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2191),
            .ce(N__2137),
            .sr(N__2087));
    defparam \generator_inst1.REGDYN7_LC_1_17_5 .C_ON=1'b0;
    defparam \generator_inst1.REGDYN7_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \generator_inst1.REGDYN7_LC_1_17_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \generator_inst1.REGDYN7_LC_1_17_5  (
            .in0(N__1570),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1536),
            .lcout(\generator_inst1.REGDYNZ0Z7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \generator_inst1.REGSTAT_83_LC_2_12_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_83_LC_2_12_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_83_LC_2_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_83_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1631),
            .lcout(\generator_inst1.REGSTATZ0Z_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2204),
            .ce(N__2147),
            .sr(N__2099));
    defparam \generator_inst1.REGSTAT_84_LC_2_12_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_84_LC_2_12_2 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_84_LC_2_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_84_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1667),
            .lcout(\generator_inst1.REGSTATZ0Z_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2204),
            .ce(N__2147),
            .sr(N__2099));
    defparam \generator_inst1.REGSTAT_81_LC_2_12_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_81_LC_2_12_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_81_LC_2_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_81_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1709),
            .lcout(\generator_inst1.REGSTATZ0Z_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2204),
            .ce(N__2147),
            .sr(N__2099));
    defparam \generator_inst1.REGSTAT_85_LC_2_12_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_85_LC_2_12_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_85_LC_2_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_85_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1661),
            .lcout(\generator_inst1.REGSTATZ0Z_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2204),
            .ce(N__2147),
            .sr(N__2099));
    defparam \generator_inst1.REGSTAT_87_LC_2_12_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_87_LC_2_12_5 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_87_LC_2_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_87_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1643),
            .lcout(\generator_inst1.REGSTATZ0Z_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2204),
            .ce(N__2147),
            .sr(N__2099));
    defparam \generator_inst1.REGSTAT_86_LC_2_12_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_86_LC_2_12_6 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_86_LC_2_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_86_LC_2_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1649),
            .lcout(\generator_inst1.REGSTATZ0Z_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2204),
            .ce(N__2147),
            .sr(N__2099));
    defparam \generator_inst1.REGSTAT_82_LC_2_12_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_82_LC_2_12_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_82_LC_2_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_82_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1637),
            .lcout(\generator_inst1.REGSTATZ0Z_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2204),
            .ce(N__2147),
            .sr(N__2099));
    defparam \generator_inst1.REGSTAT_79_LC_2_13_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_79_LC_2_13_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_79_LC_2_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_79_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1619),
            .lcout(\generator_inst1.REGSTATZ0Z_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2201),
            .ce(N__2144),
            .sr(N__2096));
    defparam \generator_inst1.REGSTAT_77_LC_2_13_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_77_LC_2_13_1 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_77_LC_2_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_77_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1703),
            .lcout(\generator_inst1.REGSTATZ0Z_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2201),
            .ce(N__2144),
            .sr(N__2096));
    defparam \generator_inst1.REGSTAT_78_LC_2_13_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_78_LC_2_13_3 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_78_LC_2_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_78_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1625),
            .lcout(\generator_inst1.REGSTATZ0Z_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2201),
            .ce(N__2144),
            .sr(N__2096));
    defparam \generator_inst1.REGSTAT_80_LC_2_13_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_80_LC_2_13_6 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_80_LC_2_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_80_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1715),
            .lcout(\generator_inst1.REGSTATZ0Z_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2201),
            .ce(N__2144),
            .sr(N__2096));
    defparam \generator_inst1.REGSTAT_15_LC_2_14_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_15_LC_2_14_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_15_LC_2_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_15_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1679),
            .lcout(\generator_inst1.REGSTATZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2197),
            .ce(N__2141),
            .sr(N__2093));
    defparam \generator_inst1.REGSTAT_76_LC_2_14_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_76_LC_2_14_2 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_76_LC_2_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_76_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1685),
            .lcout(\generator_inst1.REGSTATZ0Z_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2197),
            .ce(N__2141),
            .sr(N__2093));
    defparam \generator_inst1.REGSTAT_74_LC_2_14_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_74_LC_2_14_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_74_LC_2_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_74_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1697),
            .lcout(\generator_inst1.REGSTATZ0Z_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2197),
            .ce(N__2141),
            .sr(N__2093));
    defparam \generator_inst1.REGSTAT_73_LC_2_14_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_73_LC_2_14_5 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_73_LC_2_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_73_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1865),
            .lcout(\generator_inst1.REGSTATZ0Z_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2197),
            .ce(N__2141),
            .sr(N__2093));
    defparam \generator_inst1.REGSTAT_75_LC_2_14_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_75_LC_2_14_6 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_75_LC_2_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_75_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1691),
            .lcout(\generator_inst1.REGSTATZ0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2197),
            .ce(N__2141),
            .sr(N__2093));
    defparam \generator_inst1.REGSTAT_14_LC_2_14_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_14_LC_2_14_7 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_14_LC_2_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_14_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1838),
            .lcout(\generator_inst1.REGSTATZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2197),
            .ce(N__2141),
            .sr(N__2093));
    defparam \generator_inst1.REGSTAT_17_LC_2_15_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_17_LC_2_15_0 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_17_LC_2_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_17_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1763),
            .lcout(\generator_inst1.REGSTATZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2194),
            .ce(N__2139),
            .sr(N__2090));
    defparam \generator_inst1.REGSTAT_18_LC_2_15_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_18_LC_2_15_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_18_LC_2_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_18_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1673),
            .lcout(\generator_inst1.REGSTATZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2194),
            .ce(N__2139),
            .sr(N__2090));
    defparam \generator_inst1.REGSTAT_47_LC_2_15_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_47_LC_2_15_2 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_47_LC_2_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_47_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1991),
            .lcout(\generator_inst1.REGSTATZ0Z_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2194),
            .ce(N__2139),
            .sr(N__2090));
    defparam \generator_inst1.REGSTAT_49_LC_2_15_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_49_LC_2_15_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_49_LC_2_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_49_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1751),
            .lcout(\generator_inst1.REGSTATZ0Z_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2194),
            .ce(N__2139),
            .sr(N__2090));
    defparam \generator_inst1.REGSTAT_16_LC_2_15_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_16_LC_2_15_4 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_16_LC_2_15_4 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \generator_inst1.REGSTAT_16_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1772),
            .in3(_gnd_net_),
            .lcout(\generator_inst1.REGSTATZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2194),
            .ce(N__2139),
            .sr(N__2090));
    defparam \generator_inst1.REGSTAT_48_LC_2_15_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_48_LC_2_15_5 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_48_LC_2_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_48_LC_2_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1757),
            .lcout(\generator_inst1.REGSTATZ0Z_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2194),
            .ce(N__2139),
            .sr(N__2090));
    defparam \generator_inst1.REGSTAT_19_LC_2_15_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_19_LC_2_15_6 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_19_LC_2_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_19_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1745),
            .lcout(\generator_inst1.REGSTATZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2194),
            .ce(N__2139),
            .sr(N__2090));
    defparam \generator_inst1.REGSTAT_20_LC_2_15_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_20_LC_2_15_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_20_LC_2_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_20_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1739),
            .lcout(\generator_inst1.REGSTATZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2194),
            .ce(N__2139),
            .sr(N__2090));
    defparam \generator_inst1.REGSTAT_33_LC_2_16_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_33_LC_2_16_0 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_33_LC_2_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_33_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1814),
            .lcout(\generator_inst1.REGSTATZ0Z_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2192),
            .ce(N__2138),
            .sr(N__2086));
    defparam \generator_inst1.REGSTAT_28_LC_2_16_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_28_LC_2_16_1 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_28_LC_2_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_28_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1802),
            .lcout(\generator_inst1.REGSTATZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2192),
            .ce(N__2138),
            .sr(N__2086));
    defparam \generator_inst1.REGSTAT_29_LC_2_16_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_29_LC_2_16_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_29_LC_2_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_29_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1727),
            .lcout(\generator_inst1.REGSTATZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2192),
            .ce(N__2138),
            .sr(N__2086));
    defparam \generator_inst1.REGSTAT_30_LC_2_16_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_30_LC_2_16_4 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_30_LC_2_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_30_LC_2_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1721),
            .lcout(\generator_inst1.REGSTATZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2192),
            .ce(N__2138),
            .sr(N__2086));
    defparam \generator_inst1.REGSTAT_31_LC_2_16_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_31_LC_2_16_5 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_31_LC_2_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_31_LC_2_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1826),
            .lcout(\generator_inst1.REGSTATZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2192),
            .ce(N__2138),
            .sr(N__2086));
    defparam \generator_inst1.REGSTAT_32_LC_2_16_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_32_LC_2_16_6 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_32_LC_2_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_32_LC_2_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1820),
            .lcout(\generator_inst1.REGSTATZ0Z_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2192),
            .ce(N__2138),
            .sr(N__2086));
    defparam \generator_inst1.REGSTAT_27_LC_2_16_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_27_LC_2_16_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_27_LC_2_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_27_LC_2_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1808),
            .lcout(\generator_inst1.REGSTATZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2192),
            .ce(N__2138),
            .sr(N__2086));
    defparam \generator_inst1.REGSTAT_11_LC_3_13_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_11_LC_3_13_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_11_LC_3_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_11_LC_3_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1784),
            .lcout(\generator_inst1.REGSTATZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2205),
            .ce(N__2148),
            .sr(N__2100));
    defparam \generator_inst1.REGSTAT_12_LC_3_13_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_12_LC_3_13_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_12_LC_3_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_12_LC_3_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1796),
            .lcout(\generator_inst1.REGSTATZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2205),
            .ce(N__2148),
            .sr(N__2100));
    defparam \generator_inst1.REGSTAT_7_LC_3_13_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_7_LC_3_13_2 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_7_LC_3_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_7_LC_3_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1790),
            .lcout(\generator_inst1.REGSTATZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2205),
            .ce(N__2148),
            .sr(N__2100));
    defparam \generator_inst1.REGSTAT_6_LC_3_13_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_6_LC_3_13_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_6_LC_3_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_6_LC_3_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1973),
            .lcout(\generator_inst1.REGSTATZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2205),
            .ce(N__2148),
            .sr(N__2100));
    defparam \generator_inst1.REGSTAT_10_LC_3_13_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_10_LC_3_13_5 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_10_LC_3_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_10_LC_3_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1883),
            .lcout(\generator_inst1.REGSTATZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2205),
            .ce(N__2148),
            .sr(N__2100));
    defparam \generator_inst1.REGSTAT_8_LC_3_13_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_8_LC_3_13_6 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_8_LC_3_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_8_LC_3_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1778),
            .lcout(\generator_inst1.REGSTATZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2205),
            .ce(N__2148),
            .sr(N__2100));
    defparam \generator_inst1.REGSTAT_9_LC_3_13_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_9_LC_3_13_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_9_LC_3_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_9_LC_3_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1889),
            .lcout(\generator_inst1.REGSTATZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2205),
            .ce(N__2148),
            .sr(N__2100));
    defparam \generator_inst1.REGSTAT_62_LC_3_14_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_62_LC_3_14_0 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_62_LC_3_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_62_LC_3_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1853),
            .lcout(\generator_inst1.REGSTATZ0Z_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2202),
            .ce(N__2145),
            .sr(N__2097));
    defparam \generator_inst1.REGSTAT_64_LC_3_14_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_64_LC_3_14_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_64_LC_3_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_64_LC_3_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1871),
            .lcout(\generator_inst1.REGSTATZ0Z_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2202),
            .ce(N__2145),
            .sr(N__2097));
    defparam \generator_inst1.REGSTAT_63_LC_3_14_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_63_LC_3_14_2 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_63_LC_3_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_63_LC_3_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1877),
            .lcout(\generator_inst1.REGSTATZ0Z_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2202),
            .ce(N__2145),
            .sr(N__2097));
    defparam \generator_inst1.REGSTAT_60_LC_3_14_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_60_LC_3_14_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_60_LC_3_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_60_LC_3_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2267),
            .lcout(\generator_inst1.REGSTATZ0Z_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2202),
            .ce(N__2145),
            .sr(N__2097));
    defparam \generator_inst1.REGSTAT_72_LC_3_14_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_72_LC_3_14_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_72_LC_3_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_72_LC_3_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2039),
            .lcout(\generator_inst1.REGSTATZ0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2202),
            .ce(N__2145),
            .sr(N__2097));
    defparam \generator_inst1.REGSTAT_61_LC_3_14_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_61_LC_3_14_5 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_61_LC_3_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_61_LC_3_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1859),
            .lcout(\generator_inst1.REGSTATZ0Z_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2202),
            .ce(N__2145),
            .sr(N__2097));
    defparam \generator_inst1.REGSTAT_13_LC_3_14_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_13_LC_3_14_6 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_13_LC_3_14_6 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \generator_inst1.REGSTAT_13_LC_3_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1847),
            .in3(_gnd_net_),
            .lcout(\generator_inst1.REGSTATZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2202),
            .ce(N__2145),
            .sr(N__2097));
    defparam \generator_inst1.REGSTAT_65_LC_3_14_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_65_LC_3_14_7 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_65_LC_3_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_65_LC_3_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1832),
            .lcout(\generator_inst1.REGSTATZ0Z_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2202),
            .ce(N__2145),
            .sr(N__2097));
    defparam \generator_inst1.REGSTAT_55_LC_3_15_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_55_LC_3_15_0 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_55_LC_3_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_55_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1919),
            .lcout(\generator_inst1.REGSTATZ0Z_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2198),
            .ce(N__2142),
            .sr(N__2094));
    defparam \generator_inst1.REGSTAT_50_LC_3_15_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_50_LC_3_15_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_50_LC_3_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_50_LC_3_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1937),
            .lcout(\generator_inst1.REGSTATZ0Z_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2198),
            .ce(N__2142),
            .sr(N__2094));
    defparam \generator_inst1.REGSTAT_51_LC_3_15_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_51_LC_3_15_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_51_LC_3_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_51_LC_3_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1931),
            .lcout(\generator_inst1.REGSTATZ0Z_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2198),
            .ce(N__2142),
            .sr(N__2094));
    defparam \generator_inst1.REGSTAT_52_LC_3_15_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_52_LC_3_15_4 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_52_LC_3_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_52_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1925),
            .lcout(\generator_inst1.REGSTATZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2198),
            .ce(N__2142),
            .sr(N__2094));
    defparam \generator_inst1.REGSTAT_54_LC_3_15_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_54_LC_3_15_5 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_54_LC_3_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_54_LC_3_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1907),
            .lcout(\generator_inst1.REGSTATZ0Z_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2198),
            .ce(N__2142),
            .sr(N__2094));
    defparam \generator_inst1.REGSTAT_53_LC_3_15_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_53_LC_3_15_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_53_LC_3_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_53_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1913),
            .lcout(\generator_inst1.REGSTATZ0Z_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2198),
            .ce(N__2142),
            .sr(N__2094));
    defparam \generator_inst1.REGSTAT_43_LC_3_16_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_43_LC_3_16_1 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_43_LC_3_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_43_LC_3_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2243),
            .lcout(\generator_inst1.REGSTATZ0Z_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2195),
            .ce(N__2140),
            .sr(N__2088));
    defparam \generator_inst1.REGSTAT_44_LC_3_16_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_44_LC_3_16_2 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_44_LC_3_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_44_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1901),
            .lcout(\generator_inst1.REGSTATZ0Z_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2195),
            .ce(N__2140),
            .sr(N__2088));
    defparam \generator_inst1.REGSTAT_45_LC_3_16_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_45_LC_3_16_3 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_45_LC_3_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_45_LC_3_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1895),
            .lcout(\generator_inst1.REGSTATZ0Z_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2195),
            .ce(N__2140),
            .sr(N__2088));
    defparam \generator_inst1.REGSTAT_46_LC_3_16_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_46_LC_3_16_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_46_LC_3_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_46_LC_3_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1997),
            .lcout(\generator_inst1.REGSTATZ0Z_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2195),
            .ce(N__2140),
            .sr(N__2088));
    defparam \generator_inst1.REGSTAT_34_LC_3_16_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_34_LC_3_16_6 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_34_LC_3_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_34_LC_3_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1985),
            .lcout(\generator_inst1.REGSTATZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2195),
            .ce(N__2140),
            .sr(N__2088));
    defparam \generator_inst1.REGSTAT_0_LC_4_13_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_0_LC_4_13_1 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_0_LC_4_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_0_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\generator_inst1.REGSTATZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2207),
            .ce(N__2150),
            .sr(N__2102));
    defparam \generator_inst1.REGSTAT_2_LC_4_13_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_2_LC_4_13_2 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_2_LC_4_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_2_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1961),
            .lcout(\generator_inst1.REGSTATZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2207),
            .ce(N__2150),
            .sr(N__2102));
    defparam \generator_inst1.REGSTAT_3_LC_4_13_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_3_LC_4_13_3 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_3_LC_4_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_3_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1979),
            .lcout(\generator_inst1.REGSTATZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2207),
            .ce(N__2150),
            .sr(N__2102));
    defparam \generator_inst1.REGSTAT_5_LC_4_13_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_5_LC_4_13_4 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_5_LC_4_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_5_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1949),
            .lcout(\generator_inst1.REGSTATZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2207),
            .ce(N__2150),
            .sr(N__2102));
    defparam \generator_inst1.REGSTAT_1_LC_4_13_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_1_LC_4_13_5 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_1_LC_4_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_1_LC_4_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1967),
            .lcout(\generator_inst1.REGSTATZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2207),
            .ce(N__2150),
            .sr(N__2102));
    defparam \generator_inst1.REGSTAT_4_LC_4_13_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_4_LC_4_13_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_4_LC_4_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_4_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1955),
            .lcout(\generator_inst1.REGSTATZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2207),
            .ce(N__2150),
            .sr(N__2102));
    defparam \generator_inst1.REGSTAT_66_LC_4_14_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_66_LC_4_14_0 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_66_LC_4_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_66_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1943),
            .lcout(\generator_inst1.REGSTATZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2206),
            .ce(N__2149),
            .sr(N__2101));
    defparam \generator_inst1.REGSTAT_67_LC_4_14_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_67_LC_4_14_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_67_LC_4_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_67_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2045),
            .lcout(\generator_inst1.REGSTATZ0Z_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2206),
            .ce(N__2149),
            .sr(N__2101));
    defparam \generator_inst1.REGSTAT_69_LC_4_14_3 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_69_LC_4_14_3 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_69_LC_4_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_69_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2015),
            .lcout(\generator_inst1.REGSTATZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2206),
            .ce(N__2149),
            .sr(N__2101));
    defparam \generator_inst1.REGSTAT_71_LC_4_14_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_71_LC_4_14_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_71_LC_4_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_71_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2027),
            .lcout(\generator_inst1.REGSTATZ0Z_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2206),
            .ce(N__2149),
            .sr(N__2101));
    defparam \generator_inst1.REGSTAT_70_LC_4_14_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_70_LC_4_14_5 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_70_LC_4_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_70_LC_4_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2033),
            .lcout(\generator_inst1.REGSTATZ0Z_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2206),
            .ce(N__2149),
            .sr(N__2101));
    defparam \generator_inst1.REGSTAT_68_LC_4_14_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_68_LC_4_14_6 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_68_LC_4_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_68_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2021),
            .lcout(\generator_inst1.REGSTATZ0Z_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2206),
            .ce(N__2149),
            .sr(N__2101));
    defparam \generator_inst1.REGSTAT_56_LC_4_15_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_56_LC_4_15_0 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_56_LC_4_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_56_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2009),
            .lcout(\generator_inst1.REGSTATZ0Z_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2203),
            .ce(N__2146),
            .sr(N__2098));
    defparam \generator_inst1.REGSTAT_57_LC_4_15_1 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_57_LC_4_15_1 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_57_LC_4_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_57_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2003),
            .lcout(\generator_inst1.REGSTATZ0Z_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2203),
            .ce(N__2146),
            .sr(N__2098));
    defparam \generator_inst1.REGSTAT_36_LC_4_15_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_36_LC_4_15_2 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_36_LC_4_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_36_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2213),
            .lcout(\generator_inst1.REGSTATZ0Z_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2203),
            .ce(N__2146),
            .sr(N__2098));
    defparam \generator_inst1.REGSTAT_38_LC_4_15_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_38_LC_4_15_4 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_38_LC_4_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_38_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2255),
            .lcout(\generator_inst1.REGSTATZ0Z_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2203),
            .ce(N__2146),
            .sr(N__2098));
    defparam \generator_inst1.REGSTAT_58_LC_4_15_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_58_LC_4_15_5 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_58_LC_4_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_58_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2279),
            .lcout(\generator_inst1.REGSTATZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2203),
            .ce(N__2146),
            .sr(N__2098));
    defparam \generator_inst1.REGSTAT_59_LC_4_15_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_59_LC_4_15_6 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_59_LC_4_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_59_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2273),
            .lcout(\generator_inst1.REGSTATZ0Z_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2203),
            .ce(N__2146),
            .sr(N__2098));
    defparam \generator_inst1.REGSTAT_37_LC_4_15_7 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_37_LC_4_15_7 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_37_LC_4_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_37_LC_4_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2261),
            .lcout(\generator_inst1.REGSTATZ0Z_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2203),
            .ce(N__2146),
            .sr(N__2098));
    defparam \generator_inst1.REGSTAT_39_LC_4_16_0 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_39_LC_4_16_0 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_39_LC_4_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_39_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2249),
            .lcout(\generator_inst1.REGSTATZ0Z_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2199),
            .ce(N__2143),
            .sr(N__2091));
    defparam \generator_inst1.REGSTAT_42_LC_4_16_2 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_42_LC_4_16_2 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_42_LC_4_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_42_LC_4_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2225),
            .lcout(\generator_inst1.REGSTATZ0Z_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2199),
            .ce(N__2143),
            .sr(N__2091));
    defparam \generator_inst1.REGSTAT_40_LC_4_16_4 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_40_LC_4_16_4 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_40_LC_4_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_40_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2237),
            .lcout(\generator_inst1.REGSTATZ0Z_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2199),
            .ce(N__2143),
            .sr(N__2091));
    defparam \generator_inst1.REGSTAT_41_LC_4_16_5 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_41_LC_4_16_5 .SEQ_MODE=4'b1010;
    defparam \generator_inst1.REGSTAT_41_LC_4_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_41_LC_4_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2231),
            .lcout(\generator_inst1.REGSTATZ0Z_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2199),
            .ce(N__2143),
            .sr(N__2091));
    defparam \generator_inst1.REGSTAT_35_LC_4_16_6 .C_ON=1'b0;
    defparam \generator_inst1.REGSTAT_35_LC_4_16_6 .SEQ_MODE=4'b1011;
    defparam \generator_inst1.REGSTAT_35_LC_4_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \generator_inst1.REGSTAT_35_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2219),
            .lcout(\generator_inst1.REGSTATZ0Z_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2199),
            .ce(N__2143),
            .sr(N__2091));
endmodule // top
