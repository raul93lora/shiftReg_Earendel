-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 12 2025 16:45:17

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    signal_out : out std_logic;
    RST_N : in std_logic;
    CLK : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__1397\ : std_logic;
signal \N__1396\ : std_logic;
signal \N__1395\ : std_logic;
signal \N__1388\ : std_logic;
signal \N__1387\ : std_logic;
signal \N__1386\ : std_logic;
signal \N__1379\ : std_logic;
signal \N__1378\ : std_logic;
signal \N__1377\ : std_logic;
signal \N__1360\ : std_logic;
signal \N__1357\ : std_logic;
signal \N__1354\ : std_logic;
signal \N__1353\ : std_logic;
signal \N__1350\ : std_logic;
signal \N__1347\ : std_logic;
signal \N__1342\ : std_logic;
signal \N__1339\ : std_logic;
signal \N__1336\ : std_logic;
signal \N__1333\ : std_logic;
signal \N__1332\ : std_logic;
signal \N__1329\ : std_logic;
signal \N__1326\ : std_logic;
signal \N__1321\ : std_logic;
signal \N__1318\ : std_logic;
signal \N__1315\ : std_logic;
signal \N__1312\ : std_logic;
signal \N__1309\ : std_logic;
signal \N__1308\ : std_logic;
signal \N__1305\ : std_logic;
signal \N__1302\ : std_logic;
signal \N__1299\ : std_logic;
signal \N__1294\ : std_logic;
signal \N__1293\ : std_logic;
signal \N__1290\ : std_logic;
signal \N__1287\ : std_logic;
signal \N__1284\ : std_logic;
signal \N__1281\ : std_logic;
signal \N__1276\ : std_logic;
signal \N__1275\ : std_logic;
signal \N__1272\ : std_logic;
signal \N__1269\ : std_logic;
signal \N__1266\ : std_logic;
signal \N__1263\ : std_logic;
signal \N__1258\ : std_logic;
signal \N__1257\ : std_logic;
signal \N__1254\ : std_logic;
signal \N__1251\ : std_logic;
signal \N__1248\ : std_logic;
signal \N__1245\ : std_logic;
signal \N__1240\ : std_logic;
signal \N__1239\ : std_logic;
signal \N__1236\ : std_logic;
signal \N__1233\ : std_logic;
signal \N__1230\ : std_logic;
signal \N__1227\ : std_logic;
signal \N__1222\ : std_logic;
signal \N__1221\ : std_logic;
signal \N__1220\ : std_logic;
signal \N__1219\ : std_logic;
signal \N__1218\ : std_logic;
signal \N__1217\ : std_logic;
signal \N__1216\ : std_logic;
signal \N__1215\ : std_logic;
signal \N__1214\ : std_logic;
signal \N__1209\ : std_logic;
signal \N__1194\ : std_logic;
signal \N__1191\ : std_logic;
signal \N__1188\ : std_logic;
signal \N__1183\ : std_logic;
signal \N__1182\ : std_logic;
signal \N__1181\ : std_logic;
signal \N__1178\ : std_logic;
signal \N__1175\ : std_logic;
signal \N__1172\ : std_logic;
signal \N__1169\ : std_logic;
signal \N__1166\ : std_logic;
signal \N__1163\ : std_logic;
signal \N__1156\ : std_logic;
signal \N__1155\ : std_logic;
signal \N__1154\ : std_logic;
signal \N__1153\ : std_logic;
signal \N__1152\ : std_logic;
signal \N__1151\ : std_logic;
signal \N__1138\ : std_logic;
signal \N__1135\ : std_logic;
signal \N__1132\ : std_logic;
signal \N__1131\ : std_logic;
signal \N__1130\ : std_logic;
signal \N__1129\ : std_logic;
signal \N__1128\ : std_logic;
signal \N__1127\ : std_logic;
signal \N__1114\ : std_logic;
signal \N__1111\ : std_logic;
signal \N__1108\ : std_logic;
signal \N__1107\ : std_logic;
signal \N__1104\ : std_logic;
signal \N__1101\ : std_logic;
signal \N__1096\ : std_logic;
signal \N__1095\ : std_logic;
signal \N__1094\ : std_logic;
signal \N__1091\ : std_logic;
signal \N__1088\ : std_logic;
signal \N__1085\ : std_logic;
signal \N__1078\ : std_logic;
signal \N__1075\ : std_logic;
signal \N__1074\ : std_logic;
signal \N__1071\ : std_logic;
signal \N__1068\ : std_logic;
signal \N__1063\ : std_logic;
signal \N__1062\ : std_logic;
signal \N__1059\ : std_logic;
signal \N__1056\ : std_logic;
signal \N__1053\ : std_logic;
signal \N__1048\ : std_logic;
signal \N__1045\ : std_logic;
signal \N__1042\ : std_logic;
signal \N__1039\ : std_logic;
signal \N__1036\ : std_logic;
signal \N__1033\ : std_logic;
signal \N__1030\ : std_logic;
signal \N__1027\ : std_logic;
signal \N__1024\ : std_logic;
signal \N__1021\ : std_logic;
signal \N__1018\ : std_logic;
signal \N__1015\ : std_logic;
signal \N__1012\ : std_logic;
signal \N__1009\ : std_logic;
signal \N__1006\ : std_logic;
signal \N__1003\ : std_logic;
signal \N__1000\ : std_logic;
signal \N__999\ : std_logic;
signal \N__996\ : std_logic;
signal \N__993\ : std_logic;
signal \N__990\ : std_logic;
signal \N__987\ : std_logic;
signal \N__982\ : std_logic;
signal \N__979\ : std_logic;
signal \N__976\ : std_logic;
signal \N__973\ : std_logic;
signal \N__972\ : std_logic;
signal \N__969\ : std_logic;
signal \N__966\ : std_logic;
signal \N__961\ : std_logic;
signal \N__958\ : std_logic;
signal \N__957\ : std_logic;
signal \N__954\ : std_logic;
signal \N__951\ : std_logic;
signal \N__948\ : std_logic;
signal \N__943\ : std_logic;
signal \N__940\ : std_logic;
signal \N__937\ : std_logic;
signal \N__934\ : std_logic;
signal \N__931\ : std_logic;
signal \N__930\ : std_logic;
signal \N__927\ : std_logic;
signal \N__924\ : std_logic;
signal \N__921\ : std_logic;
signal \N__916\ : std_logic;
signal \N__913\ : std_logic;
signal \N__910\ : std_logic;
signal \N__907\ : std_logic;
signal \N__904\ : std_logic;
signal \N__903\ : std_logic;
signal \N__900\ : std_logic;
signal \N__897\ : std_logic;
signal \N__894\ : std_logic;
signal \N__891\ : std_logic;
signal \N__886\ : std_logic;
signal \N__883\ : std_logic;
signal \N__880\ : std_logic;
signal \N__877\ : std_logic;
signal \N__874\ : std_logic;
signal \N__873\ : std_logic;
signal \N__870\ : std_logic;
signal \N__867\ : std_logic;
signal \N__862\ : std_logic;
signal \N__859\ : std_logic;
signal \N__856\ : std_logic;
signal \N__855\ : std_logic;
signal \N__852\ : std_logic;
signal \N__849\ : std_logic;
signal \N__844\ : std_logic;
signal \N__841\ : std_logic;
signal \N__840\ : std_logic;
signal \N__837\ : std_logic;
signal \N__834\ : std_logic;
signal \N__829\ : std_logic;
signal \N__826\ : std_logic;
signal \N__825\ : std_logic;
signal \N__822\ : std_logic;
signal \N__819\ : std_logic;
signal \N__814\ : std_logic;
signal \N__811\ : std_logic;
signal \N__810\ : std_logic;
signal \N__807\ : std_logic;
signal \N__804\ : std_logic;
signal \N__801\ : std_logic;
signal \N__798\ : std_logic;
signal \N__793\ : std_logic;
signal \N__790\ : std_logic;
signal \N__787\ : std_logic;
signal \N__784\ : std_logic;
signal \N__781\ : std_logic;
signal \N__780\ : std_logic;
signal \N__777\ : std_logic;
signal \N__774\ : std_logic;
signal \N__769\ : std_logic;
signal \N__766\ : std_logic;
signal \N__763\ : std_logic;
signal \N__762\ : std_logic;
signal \N__759\ : std_logic;
signal \N__756\ : std_logic;
signal \N__751\ : std_logic;
signal \N__748\ : std_logic;
signal \N__745\ : std_logic;
signal \N__742\ : std_logic;
signal \N__739\ : std_logic;
signal \N__738\ : std_logic;
signal \N__737\ : std_logic;
signal \N__736\ : std_logic;
signal \N__735\ : std_logic;
signal \N__734\ : std_logic;
signal \N__733\ : std_logic;
signal \N__732\ : std_logic;
signal \N__731\ : std_logic;
signal \N__716\ : std_logic;
signal \N__711\ : std_logic;
signal \N__706\ : std_logic;
signal \N__705\ : std_logic;
signal \N__704\ : std_logic;
signal \N__703\ : std_logic;
signal \N__702\ : std_logic;
signal \N__701\ : std_logic;
signal \N__698\ : std_logic;
signal \N__697\ : std_logic;
signal \N__694\ : std_logic;
signal \N__693\ : std_logic;
signal \N__692\ : std_logic;
signal \N__689\ : std_logic;
signal \N__686\ : std_logic;
signal \N__683\ : std_logic;
signal \N__680\ : std_logic;
signal \N__677\ : std_logic;
signal \N__672\ : std_logic;
signal \N__659\ : std_logic;
signal \N__652\ : std_logic;
signal \N__651\ : std_logic;
signal \N__646\ : std_logic;
signal \N__643\ : std_logic;
signal \N__640\ : std_logic;
signal \N__637\ : std_logic;
signal \N__634\ : std_logic;
signal \N__631\ : std_logic;
signal \N__628\ : std_logic;
signal \N__625\ : std_logic;
signal \N__622\ : std_logic;
signal \N__619\ : std_logic;
signal \N__616\ : std_logic;
signal \N__613\ : std_logic;
signal \N__610\ : std_logic;
signal \N__607\ : std_logic;
signal \N__604\ : std_logic;
signal \N__601\ : std_logic;
signal \N__598\ : std_logic;
signal \N__595\ : std_logic;
signal \N__592\ : std_logic;
signal \N__589\ : std_logic;
signal \N__586\ : std_logic;
signal \N__583\ : std_logic;
signal \CLK_ibuf_gb_io_gb_input\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \generator_inst1.signal_out5_11\ : std_logic;
signal \generator_inst1.signal_out5_13_cascade_\ : std_logic;
signal \generator_inst1.signal_out5_14\ : std_logic;
signal \generator_inst1.signal_out5_15\ : std_logic;
signal \generator_inst1.signal_out5_20\ : std_logic;
signal generated_signal : std_logic;
signal signal_out_c : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_1\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_2\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_3\ : std_logic;
signal \generator_inst1.counterZ0Z_5\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_4\ : std_logic;
signal \generator_inst1.counterZ0Z_6\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_5\ : std_logic;
signal \generator_inst1.counterZ0Z_7\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_6\ : std_logic;
signal \generator_inst1.counterZ0Z_8\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_7\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_8\ : std_logic;
signal \generator_inst1.counterZ0Z_9\ : std_logic;
signal \generator_inst1.counter_RNO_0Z0Z_9\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \generator_inst1.counterZ0Z_10\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_9\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_10\ : std_logic;
signal \generator_inst1.counterZ0Z_12\ : std_logic;
signal \generator_inst1.counter_RNO_0Z0Z_12\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_11\ : std_logic;
signal \generator_inst1.counterZ0Z_13\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_12\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_13\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_14\ : std_logic;
signal \generator_inst1.counterZ0Z_16\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_15\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_16\ : std_logic;
signal \generator_inst1.counterZ0Z_17\ : std_logic;
signal \generator_inst1.counter_RNO_0Z0Z_17\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_17\ : std_logic;
signal \generator_inst1.counterZ0Z_19\ : std_logic;
signal \generator_inst1.counter_RNO_0Z0Z_19\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_18\ : std_logic;
signal \generator_inst1.counterZ0Z_20\ : std_logic;
signal \generator_inst1.counter_RNO_0Z0Z_20\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_19\ : std_logic;
signal \generator_inst1.counterZ0Z_21\ : std_logic;
signal \generator_inst1.counter_RNO_0Z0Z_21\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_20\ : std_logic;
signal \generator_inst1.counterZ0Z_22\ : std_logic;
signal \generator_inst1.counter_RNO_0Z0Z_22\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_21\ : std_logic;
signal \generator_inst1.un3_counter_1_cry_22\ : std_logic;
signal \generator_inst1.counterZ0Z_23\ : std_logic;
signal \generator_inst1.counterZ0Z_11\ : std_logic;
signal \generator_inst1.counterZ0Z_3\ : std_logic;
signal \generator_inst1.counterZ0Z_18\ : std_logic;
signal \generator_inst1.counterZ0Z_2\ : std_logic;
signal \generator_inst1.signal_out5_16\ : std_logic;
signal \generator_inst1.counterZ0Z_0\ : std_logic;
signal \CLK_c_g\ : std_logic;
signal \RST_N_c_i_g\ : std_logic;
signal \generator_inst1.counterZ0Z_4\ : std_logic;
signal \generator_inst1.counterZ0Z_1\ : std_logic;
signal \generator_inst1.counterZ0Z_14\ : std_logic;
signal \generator_inst1.counterZ0Z_15\ : std_logic;
signal \generator_inst1.signal_out5_12\ : std_logic;
signal \RST_N_c\ : std_logic;
signal \RST_N_c_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \RST_N_wire\ : std_logic;
signal signal_out_wire : std_logic;
signal \CLK_wire\ : std_logic;

begin
    \RST_N_wire\ <= RST_N;
    signal_out <= signal_out_wire;
    \CLK_wire\ <= CLK;

    \RST_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1397\,
            DIN => \N__1396\,
            DOUT => \N__1395\,
            PACKAGEPIN => \RST_N_wire\
        );

    \RST_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1397\,
            PADOUT => \N__1396\,
            PADIN => \N__1395\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RST_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \signal_out_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1388\,
            DIN => \N__1387\,
            DOUT => \N__1386\,
            PACKAGEPIN => signal_out_wire
        );

    \signal_out_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1388\,
            PADOUT => \N__1387\,
            PADIN => \N__1386\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__643\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1379\,
            DIN => \N__1378\,
            DOUT => \N__1377\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1379\,
            PADOUT => \N__1378\,
            PADIN => \N__1377\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK_ibuf_gb_io_gb_input\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__312\ : CascadeMux
    port map (
            O => \N__1360\,
            I => \N__1357\
        );

    \I__311\ : InMux
    port map (
            O => \N__1357\,
            I => \N__1354\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__1354\,
            I => \N__1350\
        );

    \I__309\ : InMux
    port map (
            O => \N__1353\,
            I => \N__1347\
        );

    \I__308\ : Odrv12
    port map (
            O => \N__1350\,
            I => \generator_inst1.counterZ0Z_21\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__1347\,
            I => \generator_inst1.counterZ0Z_21\
        );

    \I__306\ : InMux
    port map (
            O => \N__1342\,
            I => \N__1339\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__1339\,
            I => \generator_inst1.counter_RNO_0Z0Z_21\
        );

    \I__304\ : InMux
    port map (
            O => \N__1336\,
            I => \generator_inst1.un3_counter_1_cry_20\
        );

    \I__303\ : InMux
    port map (
            O => \N__1333\,
            I => \N__1329\
        );

    \I__302\ : InMux
    port map (
            O => \N__1332\,
            I => \N__1326\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__1329\,
            I => \generator_inst1.counterZ0Z_22\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__1326\,
            I => \generator_inst1.counterZ0Z_22\
        );

    \I__299\ : InMux
    port map (
            O => \N__1321\,
            I => \N__1318\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__1318\,
            I => \generator_inst1.counter_RNO_0Z0Z_22\
        );

    \I__297\ : InMux
    port map (
            O => \N__1315\,
            I => \generator_inst1.un3_counter_1_cry_21\
        );

    \I__296\ : InMux
    port map (
            O => \N__1312\,
            I => \generator_inst1.un3_counter_1_cry_22\
        );

    \I__295\ : CascadeMux
    port map (
            O => \N__1309\,
            I => \N__1305\
        );

    \I__294\ : InMux
    port map (
            O => \N__1308\,
            I => \N__1302\
        );

    \I__293\ : InMux
    port map (
            O => \N__1305\,
            I => \N__1299\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__1302\,
            I => \generator_inst1.counterZ0Z_23\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__1299\,
            I => \generator_inst1.counterZ0Z_23\
        );

    \I__290\ : InMux
    port map (
            O => \N__1294\,
            I => \N__1290\
        );

    \I__289\ : CascadeMux
    port map (
            O => \N__1293\,
            I => \N__1287\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__1290\,
            I => \N__1284\
        );

    \I__287\ : InMux
    port map (
            O => \N__1287\,
            I => \N__1281\
        );

    \I__286\ : Odrv4
    port map (
            O => \N__1284\,
            I => \generator_inst1.counterZ0Z_11\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__1281\,
            I => \generator_inst1.counterZ0Z_11\
        );

    \I__284\ : InMux
    port map (
            O => \N__1276\,
            I => \N__1272\
        );

    \I__283\ : CascadeMux
    port map (
            O => \N__1275\,
            I => \N__1269\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__1272\,
            I => \N__1266\
        );

    \I__281\ : InMux
    port map (
            O => \N__1269\,
            I => \N__1263\
        );

    \I__280\ : Odrv4
    port map (
            O => \N__1266\,
            I => \generator_inst1.counterZ0Z_3\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__1263\,
            I => \generator_inst1.counterZ0Z_3\
        );

    \I__278\ : CascadeMux
    port map (
            O => \N__1258\,
            I => \N__1254\
        );

    \I__277\ : CascadeMux
    port map (
            O => \N__1257\,
            I => \N__1251\
        );

    \I__276\ : InMux
    port map (
            O => \N__1254\,
            I => \N__1248\
        );

    \I__275\ : InMux
    port map (
            O => \N__1251\,
            I => \N__1245\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__1248\,
            I => \generator_inst1.counterZ0Z_18\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__1245\,
            I => \generator_inst1.counterZ0Z_18\
        );

    \I__272\ : InMux
    port map (
            O => \N__1240\,
            I => \N__1236\
        );

    \I__271\ : CascadeMux
    port map (
            O => \N__1239\,
            I => \N__1233\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__1236\,
            I => \N__1230\
        );

    \I__269\ : InMux
    port map (
            O => \N__1233\,
            I => \N__1227\
        );

    \I__268\ : Odrv12
    port map (
            O => \N__1230\,
            I => \generator_inst1.counterZ0Z_2\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__1227\,
            I => \generator_inst1.counterZ0Z_2\
        );

    \I__266\ : InMux
    port map (
            O => \N__1222\,
            I => \N__1209\
        );

    \I__265\ : InMux
    port map (
            O => \N__1221\,
            I => \N__1209\
        );

    \I__264\ : InMux
    port map (
            O => \N__1220\,
            I => \N__1194\
        );

    \I__263\ : InMux
    port map (
            O => \N__1219\,
            I => \N__1194\
        );

    \I__262\ : InMux
    port map (
            O => \N__1218\,
            I => \N__1194\
        );

    \I__261\ : InMux
    port map (
            O => \N__1217\,
            I => \N__1194\
        );

    \I__260\ : InMux
    port map (
            O => \N__1216\,
            I => \N__1194\
        );

    \I__259\ : InMux
    port map (
            O => \N__1215\,
            I => \N__1194\
        );

    \I__258\ : InMux
    port map (
            O => \N__1214\,
            I => \N__1194\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__1209\,
            I => \N__1191\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__1194\,
            I => \N__1188\
        );

    \I__255\ : Odrv4
    port map (
            O => \N__1191\,
            I => \generator_inst1.signal_out5_16\
        );

    \I__254\ : Odrv4
    port map (
            O => \N__1188\,
            I => \generator_inst1.signal_out5_16\
        );

    \I__253\ : CascadeMux
    port map (
            O => \N__1183\,
            I => \N__1178\
        );

    \I__252\ : InMux
    port map (
            O => \N__1182\,
            I => \N__1175\
        );

    \I__251\ : CascadeMux
    port map (
            O => \N__1181\,
            I => \N__1172\
        );

    \I__250\ : InMux
    port map (
            O => \N__1178\,
            I => \N__1169\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__1175\,
            I => \N__1166\
        );

    \I__248\ : InMux
    port map (
            O => \N__1172\,
            I => \N__1163\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__1169\,
            I => \generator_inst1.counterZ0Z_0\
        );

    \I__246\ : Odrv4
    port map (
            O => \N__1166\,
            I => \generator_inst1.counterZ0Z_0\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__1163\,
            I => \generator_inst1.counterZ0Z_0\
        );

    \I__244\ : ClkMux
    port map (
            O => \N__1156\,
            I => \N__1138\
        );

    \I__243\ : ClkMux
    port map (
            O => \N__1155\,
            I => \N__1138\
        );

    \I__242\ : ClkMux
    port map (
            O => \N__1154\,
            I => \N__1138\
        );

    \I__241\ : ClkMux
    port map (
            O => \N__1153\,
            I => \N__1138\
        );

    \I__240\ : ClkMux
    port map (
            O => \N__1152\,
            I => \N__1138\
        );

    \I__239\ : ClkMux
    port map (
            O => \N__1151\,
            I => \N__1138\
        );

    \I__238\ : GlobalMux
    port map (
            O => \N__1138\,
            I => \N__1135\
        );

    \I__237\ : gio2CtrlBuf
    port map (
            O => \N__1135\,
            I => \CLK_c_g\
        );

    \I__236\ : SRMux
    port map (
            O => \N__1132\,
            I => \N__1114\
        );

    \I__235\ : SRMux
    port map (
            O => \N__1131\,
            I => \N__1114\
        );

    \I__234\ : SRMux
    port map (
            O => \N__1130\,
            I => \N__1114\
        );

    \I__233\ : SRMux
    port map (
            O => \N__1129\,
            I => \N__1114\
        );

    \I__232\ : SRMux
    port map (
            O => \N__1128\,
            I => \N__1114\
        );

    \I__231\ : SRMux
    port map (
            O => \N__1127\,
            I => \N__1114\
        );

    \I__230\ : GlobalMux
    port map (
            O => \N__1114\,
            I => \N__1111\
        );

    \I__229\ : gio2CtrlBuf
    port map (
            O => \N__1111\,
            I => \RST_N_c_i_g\
        );

    \I__228\ : InMux
    port map (
            O => \N__1108\,
            I => \N__1104\
        );

    \I__227\ : InMux
    port map (
            O => \N__1107\,
            I => \N__1101\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__1104\,
            I => \generator_inst1.counterZ0Z_4\
        );

    \I__225\ : LocalMux
    port map (
            O => \N__1101\,
            I => \generator_inst1.counterZ0Z_4\
        );

    \I__224\ : InMux
    port map (
            O => \N__1096\,
            I => \N__1091\
        );

    \I__223\ : InMux
    port map (
            O => \N__1095\,
            I => \N__1088\
        );

    \I__222\ : InMux
    port map (
            O => \N__1094\,
            I => \N__1085\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__1091\,
            I => \generator_inst1.counterZ0Z_1\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__1088\,
            I => \generator_inst1.counterZ0Z_1\
        );

    \I__219\ : LocalMux
    port map (
            O => \N__1085\,
            I => \generator_inst1.counterZ0Z_1\
        );

    \I__218\ : CascadeMux
    port map (
            O => \N__1078\,
            I => \N__1075\
        );

    \I__217\ : InMux
    port map (
            O => \N__1075\,
            I => \N__1071\
        );

    \I__216\ : InMux
    port map (
            O => \N__1074\,
            I => \N__1068\
        );

    \I__215\ : LocalMux
    port map (
            O => \N__1071\,
            I => \generator_inst1.counterZ0Z_14\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__1068\,
            I => \generator_inst1.counterZ0Z_14\
        );

    \I__213\ : CascadeMux
    port map (
            O => \N__1063\,
            I => \N__1059\
        );

    \I__212\ : InMux
    port map (
            O => \N__1062\,
            I => \N__1056\
        );

    \I__211\ : InMux
    port map (
            O => \N__1059\,
            I => \N__1053\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__1056\,
            I => \generator_inst1.counterZ0Z_15\
        );

    \I__209\ : LocalMux
    port map (
            O => \N__1053\,
            I => \generator_inst1.counterZ0Z_15\
        );

    \I__208\ : InMux
    port map (
            O => \N__1048\,
            I => \N__1045\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__1045\,
            I => \N__1042\
        );

    \I__206\ : Odrv12
    port map (
            O => \N__1042\,
            I => \generator_inst1.signal_out5_12\
        );

    \I__205\ : InMux
    port map (
            O => \N__1039\,
            I => \N__1036\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__1036\,
            I => \N__1033\
        );

    \I__203\ : Span12Mux_v
    port map (
            O => \N__1033\,
            I => \N__1030\
        );

    \I__202\ : Odrv12
    port map (
            O => \N__1030\,
            I => \RST_N_c\
        );

    \I__201\ : IoInMux
    port map (
            O => \N__1027\,
            I => \N__1024\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__1024\,
            I => \N__1021\
        );

    \I__199\ : Span4Mux_s1_h
    port map (
            O => \N__1021\,
            I => \N__1018\
        );

    \I__198\ : Span4Mux_h
    port map (
            O => \N__1018\,
            I => \N__1015\
        );

    \I__197\ : Sp12to4
    port map (
            O => \N__1015\,
            I => \N__1012\
        );

    \I__196\ : Span12Mux_v
    port map (
            O => \N__1012\,
            I => \N__1009\
        );

    \I__195\ : Span12Mux_h
    port map (
            O => \N__1009\,
            I => \N__1006\
        );

    \I__194\ : Span12Mux_h
    port map (
            O => \N__1006\,
            I => \N__1003\
        );

    \I__193\ : Odrv12
    port map (
            O => \N__1003\,
            I => \RST_N_c_i\
        );

    \I__192\ : CascadeMux
    port map (
            O => \N__1000\,
            I => \N__996\
        );

    \I__191\ : CascadeMux
    port map (
            O => \N__999\,
            I => \N__993\
        );

    \I__190\ : InMux
    port map (
            O => \N__996\,
            I => \N__990\
        );

    \I__189\ : InMux
    port map (
            O => \N__993\,
            I => \N__987\
        );

    \I__188\ : LocalMux
    port map (
            O => \N__990\,
            I => \generator_inst1.counterZ0Z_13\
        );

    \I__187\ : LocalMux
    port map (
            O => \N__987\,
            I => \generator_inst1.counterZ0Z_13\
        );

    \I__186\ : InMux
    port map (
            O => \N__982\,
            I => \generator_inst1.un3_counter_1_cry_12\
        );

    \I__185\ : InMux
    port map (
            O => \N__979\,
            I => \generator_inst1.un3_counter_1_cry_13\
        );

    \I__184\ : InMux
    port map (
            O => \N__976\,
            I => \generator_inst1.un3_counter_1_cry_14\
        );

    \I__183\ : InMux
    port map (
            O => \N__973\,
            I => \N__969\
        );

    \I__182\ : InMux
    port map (
            O => \N__972\,
            I => \N__966\
        );

    \I__181\ : LocalMux
    port map (
            O => \N__969\,
            I => \generator_inst1.counterZ0Z_16\
        );

    \I__180\ : LocalMux
    port map (
            O => \N__966\,
            I => \generator_inst1.counterZ0Z_16\
        );

    \I__179\ : InMux
    port map (
            O => \N__961\,
            I => \generator_inst1.un3_counter_1_cry_15\
        );

    \I__178\ : InMux
    port map (
            O => \N__958\,
            I => \N__954\
        );

    \I__177\ : InMux
    port map (
            O => \N__957\,
            I => \N__951\
        );

    \I__176\ : LocalMux
    port map (
            O => \N__954\,
            I => \N__948\
        );

    \I__175\ : LocalMux
    port map (
            O => \N__951\,
            I => \generator_inst1.counterZ0Z_17\
        );

    \I__174\ : Odrv4
    port map (
            O => \N__948\,
            I => \generator_inst1.counterZ0Z_17\
        );

    \I__173\ : InMux
    port map (
            O => \N__943\,
            I => \N__940\
        );

    \I__172\ : LocalMux
    port map (
            O => \N__940\,
            I => \generator_inst1.counter_RNO_0Z0Z_17\
        );

    \I__171\ : InMux
    port map (
            O => \N__937\,
            I => \bfn_11_19_0_\
        );

    \I__170\ : InMux
    port map (
            O => \N__934\,
            I => \generator_inst1.un3_counter_1_cry_17\
        );

    \I__169\ : CascadeMux
    port map (
            O => \N__931\,
            I => \N__927\
        );

    \I__168\ : InMux
    port map (
            O => \N__930\,
            I => \N__924\
        );

    \I__167\ : InMux
    port map (
            O => \N__927\,
            I => \N__921\
        );

    \I__166\ : LocalMux
    port map (
            O => \N__924\,
            I => \generator_inst1.counterZ0Z_19\
        );

    \I__165\ : LocalMux
    port map (
            O => \N__921\,
            I => \generator_inst1.counterZ0Z_19\
        );

    \I__164\ : CascadeMux
    port map (
            O => \N__916\,
            I => \N__913\
        );

    \I__163\ : InMux
    port map (
            O => \N__913\,
            I => \N__910\
        );

    \I__162\ : LocalMux
    port map (
            O => \N__910\,
            I => \generator_inst1.counter_RNO_0Z0Z_19\
        );

    \I__161\ : InMux
    port map (
            O => \N__907\,
            I => \generator_inst1.un3_counter_1_cry_18\
        );

    \I__160\ : CascadeMux
    port map (
            O => \N__904\,
            I => \N__900\
        );

    \I__159\ : CascadeMux
    port map (
            O => \N__903\,
            I => \N__897\
        );

    \I__158\ : InMux
    port map (
            O => \N__900\,
            I => \N__894\
        );

    \I__157\ : InMux
    port map (
            O => \N__897\,
            I => \N__891\
        );

    \I__156\ : LocalMux
    port map (
            O => \N__894\,
            I => \generator_inst1.counterZ0Z_20\
        );

    \I__155\ : LocalMux
    port map (
            O => \N__891\,
            I => \generator_inst1.counterZ0Z_20\
        );

    \I__154\ : InMux
    port map (
            O => \N__886\,
            I => \N__883\
        );

    \I__153\ : LocalMux
    port map (
            O => \N__883\,
            I => \generator_inst1.counter_RNO_0Z0Z_20\
        );

    \I__152\ : InMux
    port map (
            O => \N__880\,
            I => \generator_inst1.un3_counter_1_cry_19\
        );

    \I__151\ : InMux
    port map (
            O => \N__877\,
            I => \generator_inst1.un3_counter_1_cry_3\
        );

    \I__150\ : InMux
    port map (
            O => \N__874\,
            I => \N__870\
        );

    \I__149\ : InMux
    port map (
            O => \N__873\,
            I => \N__867\
        );

    \I__148\ : LocalMux
    port map (
            O => \N__870\,
            I => \generator_inst1.counterZ0Z_5\
        );

    \I__147\ : LocalMux
    port map (
            O => \N__867\,
            I => \generator_inst1.counterZ0Z_5\
        );

    \I__146\ : InMux
    port map (
            O => \N__862\,
            I => \generator_inst1.un3_counter_1_cry_4\
        );

    \I__145\ : InMux
    port map (
            O => \N__859\,
            I => \N__856\
        );

    \I__144\ : LocalMux
    port map (
            O => \N__856\,
            I => \N__852\
        );

    \I__143\ : InMux
    port map (
            O => \N__855\,
            I => \N__849\
        );

    \I__142\ : Odrv4
    port map (
            O => \N__852\,
            I => \generator_inst1.counterZ0Z_6\
        );

    \I__141\ : LocalMux
    port map (
            O => \N__849\,
            I => \generator_inst1.counterZ0Z_6\
        );

    \I__140\ : InMux
    port map (
            O => \N__844\,
            I => \generator_inst1.un3_counter_1_cry_5\
        );

    \I__139\ : InMux
    port map (
            O => \N__841\,
            I => \N__837\
        );

    \I__138\ : InMux
    port map (
            O => \N__840\,
            I => \N__834\
        );

    \I__137\ : LocalMux
    port map (
            O => \N__837\,
            I => \generator_inst1.counterZ0Z_7\
        );

    \I__136\ : LocalMux
    port map (
            O => \N__834\,
            I => \generator_inst1.counterZ0Z_7\
        );

    \I__135\ : InMux
    port map (
            O => \N__829\,
            I => \generator_inst1.un3_counter_1_cry_6\
        );

    \I__134\ : InMux
    port map (
            O => \N__826\,
            I => \N__822\
        );

    \I__133\ : InMux
    port map (
            O => \N__825\,
            I => \N__819\
        );

    \I__132\ : LocalMux
    port map (
            O => \N__822\,
            I => \generator_inst1.counterZ0Z_8\
        );

    \I__131\ : LocalMux
    port map (
            O => \N__819\,
            I => \generator_inst1.counterZ0Z_8\
        );

    \I__130\ : InMux
    port map (
            O => \N__814\,
            I => \generator_inst1.un3_counter_1_cry_7\
        );

    \I__129\ : InMux
    port map (
            O => \N__811\,
            I => \N__807\
        );

    \I__128\ : CascadeMux
    port map (
            O => \N__810\,
            I => \N__804\
        );

    \I__127\ : LocalMux
    port map (
            O => \N__807\,
            I => \N__801\
        );

    \I__126\ : InMux
    port map (
            O => \N__804\,
            I => \N__798\
        );

    \I__125\ : Odrv4
    port map (
            O => \N__801\,
            I => \generator_inst1.counterZ0Z_9\
        );

    \I__124\ : LocalMux
    port map (
            O => \N__798\,
            I => \generator_inst1.counterZ0Z_9\
        );

    \I__123\ : InMux
    port map (
            O => \N__793\,
            I => \N__790\
        );

    \I__122\ : LocalMux
    port map (
            O => \N__790\,
            I => \generator_inst1.counter_RNO_0Z0Z_9\
        );

    \I__121\ : InMux
    port map (
            O => \N__787\,
            I => \bfn_11_18_0_\
        );

    \I__120\ : InMux
    port map (
            O => \N__784\,
            I => \N__781\
        );

    \I__119\ : LocalMux
    port map (
            O => \N__781\,
            I => \N__777\
        );

    \I__118\ : InMux
    port map (
            O => \N__780\,
            I => \N__774\
        );

    \I__117\ : Odrv4
    port map (
            O => \N__777\,
            I => \generator_inst1.counterZ0Z_10\
        );

    \I__116\ : LocalMux
    port map (
            O => \N__774\,
            I => \generator_inst1.counterZ0Z_10\
        );

    \I__115\ : InMux
    port map (
            O => \N__769\,
            I => \generator_inst1.un3_counter_1_cry_9\
        );

    \I__114\ : InMux
    port map (
            O => \N__766\,
            I => \generator_inst1.un3_counter_1_cry_10\
        );

    \I__113\ : InMux
    port map (
            O => \N__763\,
            I => \N__759\
        );

    \I__112\ : InMux
    port map (
            O => \N__762\,
            I => \N__756\
        );

    \I__111\ : LocalMux
    port map (
            O => \N__759\,
            I => \generator_inst1.counterZ0Z_12\
        );

    \I__110\ : LocalMux
    port map (
            O => \N__756\,
            I => \generator_inst1.counterZ0Z_12\
        );

    \I__109\ : CascadeMux
    port map (
            O => \N__751\,
            I => \N__748\
        );

    \I__108\ : InMux
    port map (
            O => \N__748\,
            I => \N__745\
        );

    \I__107\ : LocalMux
    port map (
            O => \N__745\,
            I => \generator_inst1.counter_RNO_0Z0Z_12\
        );

    \I__106\ : InMux
    port map (
            O => \N__742\,
            I => \generator_inst1.un3_counter_1_cry_11\
        );

    \I__105\ : InMux
    port map (
            O => \N__739\,
            I => \N__716\
        );

    \I__104\ : InMux
    port map (
            O => \N__738\,
            I => \N__716\
        );

    \I__103\ : InMux
    port map (
            O => \N__737\,
            I => \N__716\
        );

    \I__102\ : InMux
    port map (
            O => \N__736\,
            I => \N__716\
        );

    \I__101\ : InMux
    port map (
            O => \N__735\,
            I => \N__716\
        );

    \I__100\ : InMux
    port map (
            O => \N__734\,
            I => \N__716\
        );

    \I__99\ : InMux
    port map (
            O => \N__733\,
            I => \N__716\
        );

    \I__98\ : InMux
    port map (
            O => \N__732\,
            I => \N__711\
        );

    \I__97\ : InMux
    port map (
            O => \N__731\,
            I => \N__711\
        );

    \I__96\ : LocalMux
    port map (
            O => \N__716\,
            I => \generator_inst1.signal_out5_15\
        );

    \I__95\ : LocalMux
    port map (
            O => \N__711\,
            I => \generator_inst1.signal_out5_15\
        );

    \I__94\ : CascadeMux
    port map (
            O => \N__706\,
            I => \N__698\
        );

    \I__93\ : CascadeMux
    port map (
            O => \N__705\,
            I => \N__694\
        );

    \I__92\ : CascadeMux
    port map (
            O => \N__704\,
            I => \N__689\
        );

    \I__91\ : CascadeMux
    port map (
            O => \N__703\,
            I => \N__686\
        );

    \I__90\ : CascadeMux
    port map (
            O => \N__702\,
            I => \N__683\
        );

    \I__89\ : CascadeMux
    port map (
            O => \N__701\,
            I => \N__680\
        );

    \I__88\ : InMux
    port map (
            O => \N__698\,
            I => \N__677\
        );

    \I__87\ : InMux
    port map (
            O => \N__697\,
            I => \N__672\
        );

    \I__86\ : InMux
    port map (
            O => \N__694\,
            I => \N__672\
        );

    \I__85\ : InMux
    port map (
            O => \N__693\,
            I => \N__659\
        );

    \I__84\ : InMux
    port map (
            O => \N__692\,
            I => \N__659\
        );

    \I__83\ : InMux
    port map (
            O => \N__689\,
            I => \N__659\
        );

    \I__82\ : InMux
    port map (
            O => \N__686\,
            I => \N__659\
        );

    \I__81\ : InMux
    port map (
            O => \N__683\,
            I => \N__659\
        );

    \I__80\ : InMux
    port map (
            O => \N__680\,
            I => \N__659\
        );

    \I__79\ : LocalMux
    port map (
            O => \N__677\,
            I => \generator_inst1.signal_out5_20\
        );

    \I__78\ : LocalMux
    port map (
            O => \N__672\,
            I => \generator_inst1.signal_out5_20\
        );

    \I__77\ : LocalMux
    port map (
            O => \N__659\,
            I => \generator_inst1.signal_out5_20\
        );

    \I__76\ : InMux
    port map (
            O => \N__652\,
            I => \N__646\
        );

    \I__75\ : InMux
    port map (
            O => \N__651\,
            I => \N__646\
        );

    \I__74\ : LocalMux
    port map (
            O => \N__646\,
            I => generated_signal
        );

    \I__73\ : IoInMux
    port map (
            O => \N__643\,
            I => \N__640\
        );

    \I__72\ : LocalMux
    port map (
            O => \N__640\,
            I => \N__637\
        );

    \I__71\ : IoSpan4Mux
    port map (
            O => \N__637\,
            I => \N__634\
        );

    \I__70\ : Span4Mux_s2_v
    port map (
            O => \N__634\,
            I => \N__631\
        );

    \I__69\ : Sp12to4
    port map (
            O => \N__631\,
            I => \N__628\
        );

    \I__68\ : Span12Mux_v
    port map (
            O => \N__628\,
            I => \N__625\
        );

    \I__67\ : Span12Mux_h
    port map (
            O => \N__625\,
            I => \N__622\
        );

    \I__66\ : Odrv12
    port map (
            O => \N__622\,
            I => signal_out_c
        );

    \I__65\ : InMux
    port map (
            O => \N__619\,
            I => \generator_inst1.un3_counter_1_cry_1\
        );

    \I__64\ : InMux
    port map (
            O => \N__616\,
            I => \generator_inst1.un3_counter_1_cry_2\
        );

    \I__63\ : InMux
    port map (
            O => \N__613\,
            I => \N__610\
        );

    \I__62\ : LocalMux
    port map (
            O => \N__610\,
            I => \generator_inst1.signal_out5_11\
        );

    \I__61\ : CascadeMux
    port map (
            O => \N__607\,
            I => \generator_inst1.signal_out5_13_cascade_\
        );

    \I__60\ : InMux
    port map (
            O => \N__604\,
            I => \N__601\
        );

    \I__59\ : LocalMux
    port map (
            O => \N__601\,
            I => \generator_inst1.signal_out5_14\
        );

    \I__58\ : IoInMux
    port map (
            O => \N__598\,
            I => \N__595\
        );

    \I__57\ : LocalMux
    port map (
            O => \N__595\,
            I => \N__592\
        );

    \I__56\ : IoSpan4Mux
    port map (
            O => \N__592\,
            I => \N__589\
        );

    \I__55\ : IoSpan4Mux
    port map (
            O => \N__589\,
            I => \N__586\
        );

    \I__54\ : IoSpan4Mux
    port map (
            O => \N__586\,
            I => \N__583\
        );

    \I__53\ : Odrv4
    port map (
            O => \N__583\,
            I => \CLK_ibuf_gb_io_gb_input\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \generator_inst1.un3_counter_1_cry_8\,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \generator_inst1.un3_counter_1_cry_16\,
            carryinitout => \bfn_11_19_0_\
        );

    \CLK_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__598\,
            GLOBALBUFFEROUTPUT => \CLK_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \RST_N_ibuf_RNIBJGC_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__1027\,
            GLOBALBUFFEROUTPUT => \RST_N_c_i_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \generator_inst1.counter_0_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__1221\,
            in1 => \N__731\,
            in2 => \N__1183\,
            in3 => \N__697\,
            lcout => \generator_inst1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1151\,
            ce => 'H',
            sr => \N__1127\
        );

    \generator_inst1.counter_9_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__732\,
            in1 => \N__1222\,
            in2 => \N__705\,
            in3 => \N__793\,
            lcout => \generator_inst1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1151\,
            ce => 'H',
            sr => \N__1127\
        );

    \generator_inst1.counter_RNI30RL1_12_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__958\,
            in1 => \N__763\,
            in2 => \N__904\,
            in3 => \N__930\,
            lcout => \generator_inst1.signal_out5_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.counter_RNIIF331_23_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000001"
        )
    port map (
            in0 => \N__973\,
            in1 => \N__874\,
            in2 => \N__1309\,
            in3 => \_gnd_net_\,
            lcout => \generator_inst1.signal_out5_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.counter_RNIM0V51_6_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__811\,
            in1 => \N__841\,
            in2 => \N__1000\,
            in3 => \N__859\,
            lcout => \generator_inst1.signal_out5_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.counter_RNICPIG1_8_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__784\,
            in1 => \N__826\,
            in2 => \N__1360\,
            in3 => \N__1332\,
            lcout => OPEN,
            ltout => \generator_inst1.signal_out5_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.counter_RNITVOK5_1_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__613\,
            in1 => \N__1048\,
            in2 => \N__607\,
            in3 => \N__604\,
            lcout => \generator_inst1.signal_out5_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.signal_out_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__739\,
            in1 => \N__651\,
            in2 => \N__704\,
            in3 => \N__1220\,
            lcout => generated_signal,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1154\,
            ce => 'H',
            sr => \N__1129\
        );

    \generator_inst1.counter_21_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__1218\,
            in1 => \N__737\,
            in2 => \N__706\,
            in3 => \N__1342\,
            lcout => \generator_inst1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1154\,
            ce => 'H',
            sr => \N__1129\
        );

    \generator_inst1.counter_22_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__738\,
            in1 => \N__1219\,
            in2 => \N__703\,
            in3 => \N__1321\,
            lcout => \generator_inst1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1154\,
            ce => 'H',
            sr => \N__1129\
        );

    \generator_inst1.counter_12_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__1214\,
            in1 => \N__733\,
            in2 => \N__751\,
            in3 => \N__692\,
            lcout => \generator_inst1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1154\,
            ce => 'H',
            sr => \N__1129\
        );

    \generator_inst1.counter_17_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__734\,
            in1 => \N__1215\,
            in2 => \N__701\,
            in3 => \N__943\,
            lcout => \generator_inst1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1154\,
            ce => 'H',
            sr => \N__1129\
        );

    \generator_inst1.counter_19_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__1216\,
            in1 => \N__735\,
            in2 => \N__916\,
            in3 => \N__693\,
            lcout => \generator_inst1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1154\,
            ce => 'H',
            sr => \N__1129\
        );

    \generator_inst1.counter_20_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__736\,
            in1 => \N__1217\,
            in2 => \N__702\,
            in3 => \N__886\,
            lcout => \generator_inst1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1154\,
            ce => 'H',
            sr => \N__1129\
        );

    \receptor_inst1.signal_out_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__652\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => signal_out_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1154\,
            ce => 'H',
            sr => \N__1129\
        );

    \generator_inst1.un3_counter_1_cry_1_c_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1094\,
            in2 => \N__1181\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \generator_inst1.un3_counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.counter_2_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1239\,
            in3 => \N__619\,
            lcout => \generator_inst1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_1\,
            carryout => \generator_inst1.un3_counter_1_cry_2\,
            clk => \N__1152\,
            ce => 'H',
            sr => \N__1128\
        );

    \generator_inst1.counter_3_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1275\,
            in3 => \N__616\,
            lcout => \generator_inst1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_2\,
            carryout => \generator_inst1.un3_counter_1_cry_3\,
            clk => \N__1152\,
            ce => 'H',
            sr => \N__1128\
        );

    \generator_inst1.counter_4_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1107\,
            in2 => \_gnd_net_\,
            in3 => \N__877\,
            lcout => \generator_inst1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_3\,
            carryout => \generator_inst1.un3_counter_1_cry_4\,
            clk => \N__1152\,
            ce => 'H',
            sr => \N__1128\
        );

    \generator_inst1.counter_5_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__873\,
            in2 => \_gnd_net_\,
            in3 => \N__862\,
            lcout => \generator_inst1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_4\,
            carryout => \generator_inst1.un3_counter_1_cry_5\,
            clk => \N__1152\,
            ce => 'H',
            sr => \N__1128\
        );

    \generator_inst1.counter_6_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__855\,
            in2 => \_gnd_net_\,
            in3 => \N__844\,
            lcout => \generator_inst1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_5\,
            carryout => \generator_inst1.un3_counter_1_cry_6\,
            clk => \N__1152\,
            ce => 'H',
            sr => \N__1128\
        );

    \generator_inst1.counter_7_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__840\,
            in2 => \_gnd_net_\,
            in3 => \N__829\,
            lcout => \generator_inst1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_6\,
            carryout => \generator_inst1.un3_counter_1_cry_7\,
            clk => \N__1152\,
            ce => 'H',
            sr => \N__1128\
        );

    \generator_inst1.counter_8_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__825\,
            in2 => \_gnd_net_\,
            in3 => \N__814\,
            lcout => \generator_inst1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_7\,
            carryout => \generator_inst1.un3_counter_1_cry_8\,
            clk => \N__1152\,
            ce => 'H',
            sr => \N__1128\
        );

    \generator_inst1.counter_RNO_0_9_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__810\,
            in3 => \N__787\,
            lcout => \generator_inst1.counter_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \generator_inst1.un3_counter_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.counter_10_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__780\,
            in2 => \_gnd_net_\,
            in3 => \N__769\,
            lcout => \generator_inst1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_9\,
            carryout => \generator_inst1.un3_counter_1_cry_10\,
            clk => \N__1155\,
            ce => 'H',
            sr => \N__1130\
        );

    \generator_inst1.counter_11_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1293\,
            in3 => \N__766\,
            lcout => \generator_inst1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_10\,
            carryout => \generator_inst1.un3_counter_1_cry_11\,
            clk => \N__1155\,
            ce => 'H',
            sr => \N__1130\
        );

    \generator_inst1.counter_RNO_0_12_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__762\,
            in2 => \_gnd_net_\,
            in3 => \N__742\,
            lcout => \generator_inst1.counter_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_11\,
            carryout => \generator_inst1.un3_counter_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.counter_13_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__999\,
            in3 => \N__982\,
            lcout => \generator_inst1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_12\,
            carryout => \generator_inst1.un3_counter_1_cry_13\,
            clk => \N__1155\,
            ce => 'H',
            sr => \N__1130\
        );

    \generator_inst1.counter_14_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1074\,
            in2 => \_gnd_net_\,
            in3 => \N__979\,
            lcout => \generator_inst1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_13\,
            carryout => \generator_inst1.un3_counter_1_cry_14\,
            clk => \N__1155\,
            ce => 'H',
            sr => \N__1130\
        );

    \generator_inst1.counter_15_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1063\,
            in3 => \N__976\,
            lcout => \generator_inst1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_14\,
            carryout => \generator_inst1.un3_counter_1_cry_15\,
            clk => \N__1155\,
            ce => 'H',
            sr => \N__1130\
        );

    \generator_inst1.counter_16_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__972\,
            in2 => \_gnd_net_\,
            in3 => \N__961\,
            lcout => \generator_inst1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_15\,
            carryout => \generator_inst1.un3_counter_1_cry_16\,
            clk => \N__1155\,
            ce => 'H',
            sr => \N__1130\
        );

    \generator_inst1.counter_RNO_0_17_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__957\,
            in2 => \_gnd_net_\,
            in3 => \N__937\,
            lcout => \generator_inst1.counter_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \generator_inst1.un3_counter_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.counter_18_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1257\,
            in3 => \N__934\,
            lcout => \generator_inst1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_17\,
            carryout => \generator_inst1.un3_counter_1_cry_18\,
            clk => \N__1156\,
            ce => 'H',
            sr => \N__1132\
        );

    \generator_inst1.counter_RNO_0_19_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__931\,
            in3 => \N__907\,
            lcout => \generator_inst1.counter_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_18\,
            carryout => \generator_inst1.un3_counter_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.counter_RNO_0_20_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__903\,
            in3 => \N__880\,
            lcout => \generator_inst1.counter_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_19\,
            carryout => \generator_inst1.un3_counter_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.counter_RNO_0_21_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1353\,
            in2 => \_gnd_net_\,
            in3 => \N__1336\,
            lcout => \generator_inst1.counter_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_20\,
            carryout => \generator_inst1.un3_counter_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.counter_RNO_0_22_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1333\,
            in2 => \_gnd_net_\,
            in3 => \N__1315\,
            lcout => \generator_inst1.counter_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \generator_inst1.un3_counter_1_cry_21\,
            carryout => \generator_inst1.un3_counter_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.counter_23_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1308\,
            in2 => \_gnd_net_\,
            in3 => \N__1312\,
            lcout => \generator_inst1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1156\,
            ce => 'H',
            sr => \N__1132\
        );

    \generator_inst1.counter_RNISM7B1_2_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1294\,
            in1 => \N__1276\,
            in2 => \N__1258\,
            in3 => \N__1240\,
            lcout => \generator_inst1.signal_out5_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.counter_1_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1182\,
            in2 => \_gnd_net_\,
            in3 => \N__1096\,
            lcout => \generator_inst1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1153\,
            ce => 'H',
            sr => \N__1131\
        );

    \generator_inst1.counter_RNISM7B1_1_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1108\,
            in1 => \N__1095\,
            in2 => \N__1078\,
            in3 => \N__1062\,
            lcout => \generator_inst1.signal_out5_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RST_N_ibuf_RNIBJGC_LC_30_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1039\,
            lcout => \RST_N_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
