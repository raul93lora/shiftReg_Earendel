-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 13 2025 09:41:53

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    signal_out : out std_logic;
    CLK : in std_logic;
    SELSTAT : in std_logic;
    SELDYN : in std_logic;
    RST_N : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__2336\ : std_logic;
signal \N__2335\ : std_logic;
signal \N__2334\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2323\ : std_logic;
signal \N__2316\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2314\ : std_logic;
signal \N__2307\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2296\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2273\ : std_logic;
signal \N__2270\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2252\ : std_logic;
signal \N__2249\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2240\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2225\ : std_logic;
signal \N__2222\ : std_logic;
signal \N__2219\ : std_logic;
signal \N__2216\ : std_logic;
signal \N__2213\ : std_logic;
signal \N__2210\ : std_logic;
signal \N__2207\ : std_logic;
signal \N__2206\ : std_logic;
signal \N__2205\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2203\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2200\ : std_logic;
signal \N__2199\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2197\ : std_logic;
signal \N__2196\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2194\ : std_logic;
signal \N__2193\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2191\ : std_logic;
signal \N__2156\ : std_logic;
signal \N__2153\ : std_logic;
signal \N__2150\ : std_logic;
signal \N__2149\ : std_logic;
signal \N__2148\ : std_logic;
signal \N__2147\ : std_logic;
signal \N__2146\ : std_logic;
signal \N__2145\ : std_logic;
signal \N__2144\ : std_logic;
signal \N__2143\ : std_logic;
signal \N__2142\ : std_logic;
signal \N__2141\ : std_logic;
signal \N__2140\ : std_logic;
signal \N__2139\ : std_logic;
signal \N__2138\ : std_logic;
signal \N__2137\ : std_logic;
signal \N__2108\ : std_logic;
signal \N__2105\ : std_logic;
signal \N__2102\ : std_logic;
signal \N__2101\ : std_logic;
signal \N__2100\ : std_logic;
signal \N__2099\ : std_logic;
signal \N__2098\ : std_logic;
signal \N__2097\ : std_logic;
signal \N__2096\ : std_logic;
signal \N__2095\ : std_logic;
signal \N__2094\ : std_logic;
signal \N__2093\ : std_logic;
signal \N__2092\ : std_logic;
signal \N__2091\ : std_logic;
signal \N__2090\ : std_logic;
signal \N__2089\ : std_logic;
signal \N__2088\ : std_logic;
signal \N__2087\ : std_logic;
signal \N__2086\ : std_logic;
signal \N__2051\ : std_logic;
signal \N__2048\ : std_logic;
signal \N__2045\ : std_logic;
signal \N__2042\ : std_logic;
signal \N__2039\ : std_logic;
signal \N__2036\ : std_logic;
signal \N__2033\ : std_logic;
signal \N__2030\ : std_logic;
signal \N__2027\ : std_logic;
signal \N__2024\ : std_logic;
signal \N__2021\ : std_logic;
signal \N__2018\ : std_logic;
signal \N__2015\ : std_logic;
signal \N__2012\ : std_logic;
signal \N__2009\ : std_logic;
signal \N__2006\ : std_logic;
signal \N__2003\ : std_logic;
signal \N__2000\ : std_logic;
signal \N__1997\ : std_logic;
signal \N__1994\ : std_logic;
signal \N__1991\ : std_logic;
signal \N__1988\ : std_logic;
signal \N__1985\ : std_logic;
signal \N__1982\ : std_logic;
signal \N__1979\ : std_logic;
signal \N__1976\ : std_logic;
signal \N__1973\ : std_logic;
signal \N__1970\ : std_logic;
signal \N__1967\ : std_logic;
signal \N__1964\ : std_logic;
signal \N__1961\ : std_logic;
signal \N__1958\ : std_logic;
signal \N__1955\ : std_logic;
signal \N__1952\ : std_logic;
signal \N__1949\ : std_logic;
signal \N__1946\ : std_logic;
signal \N__1943\ : std_logic;
signal \N__1940\ : std_logic;
signal \N__1937\ : std_logic;
signal \N__1934\ : std_logic;
signal \N__1931\ : std_logic;
signal \N__1928\ : std_logic;
signal \N__1925\ : std_logic;
signal \N__1922\ : std_logic;
signal \N__1919\ : std_logic;
signal \N__1916\ : std_logic;
signal \N__1913\ : std_logic;
signal \N__1910\ : std_logic;
signal \N__1907\ : std_logic;
signal \N__1904\ : std_logic;
signal \N__1901\ : std_logic;
signal \N__1898\ : std_logic;
signal \N__1895\ : std_logic;
signal \N__1892\ : std_logic;
signal \N__1889\ : std_logic;
signal \N__1886\ : std_logic;
signal \N__1883\ : std_logic;
signal \N__1880\ : std_logic;
signal \N__1877\ : std_logic;
signal \N__1874\ : std_logic;
signal \N__1871\ : std_logic;
signal \N__1868\ : std_logic;
signal \N__1865\ : std_logic;
signal \N__1862\ : std_logic;
signal \N__1859\ : std_logic;
signal \N__1856\ : std_logic;
signal \N__1853\ : std_logic;
signal \N__1850\ : std_logic;
signal \N__1847\ : std_logic;
signal \N__1844\ : std_logic;
signal \N__1841\ : std_logic;
signal \N__1838\ : std_logic;
signal \N__1835\ : std_logic;
signal \N__1832\ : std_logic;
signal \N__1829\ : std_logic;
signal \N__1826\ : std_logic;
signal \N__1823\ : std_logic;
signal \N__1820\ : std_logic;
signal \N__1817\ : std_logic;
signal \N__1814\ : std_logic;
signal \N__1811\ : std_logic;
signal \N__1808\ : std_logic;
signal \N__1805\ : std_logic;
signal \N__1802\ : std_logic;
signal \N__1799\ : std_logic;
signal \N__1796\ : std_logic;
signal \N__1793\ : std_logic;
signal \N__1790\ : std_logic;
signal \N__1787\ : std_logic;
signal \N__1784\ : std_logic;
signal \N__1781\ : std_logic;
signal \N__1778\ : std_logic;
signal \N__1775\ : std_logic;
signal \N__1772\ : std_logic;
signal \N__1769\ : std_logic;
signal \N__1766\ : std_logic;
signal \N__1763\ : std_logic;
signal \N__1760\ : std_logic;
signal \N__1757\ : std_logic;
signal \N__1754\ : std_logic;
signal \N__1751\ : std_logic;
signal \N__1748\ : std_logic;
signal \N__1745\ : std_logic;
signal \N__1742\ : std_logic;
signal \N__1739\ : std_logic;
signal \N__1736\ : std_logic;
signal \N__1733\ : std_logic;
signal \N__1730\ : std_logic;
signal \N__1727\ : std_logic;
signal \N__1724\ : std_logic;
signal \N__1721\ : std_logic;
signal \N__1718\ : std_logic;
signal \N__1715\ : std_logic;
signal \N__1712\ : std_logic;
signal \N__1709\ : std_logic;
signal \N__1706\ : std_logic;
signal \N__1703\ : std_logic;
signal \N__1700\ : std_logic;
signal \N__1697\ : std_logic;
signal \N__1694\ : std_logic;
signal \N__1691\ : std_logic;
signal \N__1688\ : std_logic;
signal \N__1685\ : std_logic;
signal \N__1682\ : std_logic;
signal \N__1679\ : std_logic;
signal \N__1676\ : std_logic;
signal \N__1673\ : std_logic;
signal \N__1670\ : std_logic;
signal \N__1667\ : std_logic;
signal \N__1664\ : std_logic;
signal \N__1661\ : std_logic;
signal \N__1658\ : std_logic;
signal \N__1655\ : std_logic;
signal \N__1652\ : std_logic;
signal \N__1649\ : std_logic;
signal \N__1646\ : std_logic;
signal \N__1643\ : std_logic;
signal \N__1640\ : std_logic;
signal \N__1637\ : std_logic;
signal \N__1634\ : std_logic;
signal \N__1631\ : std_logic;
signal \N__1628\ : std_logic;
signal \N__1625\ : std_logic;
signal \N__1622\ : std_logic;
signal \N__1619\ : std_logic;
signal \N__1616\ : std_logic;
signal \N__1613\ : std_logic;
signal \N__1610\ : std_logic;
signal \N__1607\ : std_logic;
signal \N__1604\ : std_logic;
signal \N__1601\ : std_logic;
signal \N__1598\ : std_logic;
signal \N__1595\ : std_logic;
signal \N__1592\ : std_logic;
signal \N__1589\ : std_logic;
signal \N__1586\ : std_logic;
signal \N__1583\ : std_logic;
signal \N__1580\ : std_logic;
signal \N__1577\ : std_logic;
signal \N__1574\ : std_logic;
signal \N__1571\ : std_logic;
signal \N__1570\ : std_logic;
signal \N__1567\ : std_logic;
signal \N__1564\ : std_logic;
signal \N__1559\ : std_logic;
signal \N__1556\ : std_logic;
signal \N__1555\ : std_logic;
signal \N__1552\ : std_logic;
signal \N__1549\ : std_logic;
signal \N__1544\ : std_logic;
signal \N__1543\ : std_logic;
signal \N__1540\ : std_logic;
signal \N__1537\ : std_logic;
signal \N__1536\ : std_logic;
signal \N__1531\ : std_logic;
signal \N__1528\ : std_logic;
signal \N__1523\ : std_logic;
signal \N__1520\ : std_logic;
signal \N__1517\ : std_logic;
signal \N__1514\ : std_logic;
signal \N__1511\ : std_logic;
signal \N__1508\ : std_logic;
signal \N__1505\ : std_logic;
signal \N__1502\ : std_logic;
signal \N__1499\ : std_logic;
signal \N__1496\ : std_logic;
signal \N__1493\ : std_logic;
signal \N__1490\ : std_logic;
signal \N__1487\ : std_logic;
signal \N__1484\ : std_logic;
signal \N__1481\ : std_logic;
signal \N__1478\ : std_logic;
signal \N__1475\ : std_logic;
signal \N__1472\ : std_logic;
signal \N__1469\ : std_logic;
signal \N__1466\ : std_logic;
signal \N__1463\ : std_logic;
signal \N__1460\ : std_logic;
signal \N__1457\ : std_logic;
signal \N__1454\ : std_logic;
signal \N__1451\ : std_logic;
signal \N__1448\ : std_logic;
signal \N__1445\ : std_logic;
signal \N__1442\ : std_logic;
signal \N__1439\ : std_logic;
signal \N__1436\ : std_logic;
signal \N__1433\ : std_logic;
signal \N__1430\ : std_logic;
signal \N__1427\ : std_logic;
signal \N__1424\ : std_logic;
signal \N__1421\ : std_logic;
signal \N__1418\ : std_logic;
signal \N__1415\ : std_logic;
signal \N__1412\ : std_logic;
signal \N__1409\ : std_logic;
signal \N__1406\ : std_logic;
signal \N__1403\ : std_logic;
signal \N__1400\ : std_logic;
signal \N__1397\ : std_logic;
signal \N__1394\ : std_logic;
signal \N__1391\ : std_logic;
signal \N__1388\ : std_logic;
signal \N__1385\ : std_logic;
signal \N__1382\ : std_logic;
signal \N__1379\ : std_logic;
signal \N__1376\ : std_logic;
signal \N__1373\ : std_logic;
signal \N__1370\ : std_logic;
signal \VCCG0\ : std_logic;
signal \RST_N_c\ : std_logic;
signal \RST_N_c_i\ : std_logic;
signal generated_signal : std_logic;
signal signal_out_c : std_logic;
signal \generator_inst1.REGDYNZ0Z_8\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_12\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_13\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_14\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_15\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_11\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_9\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_10\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_1\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_2\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_6\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_7\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_5\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_3\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_4\ : std_logic;
signal \generator_inst1.REGDYNZ0Z_0\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_24\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_25\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_22\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_23\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_21\ : std_logic;
signal \SELSTAT_c\ : std_logic;
signal \SELDYN_c\ : std_logic;
signal \generator_inst1.REGDYNZ0Z7\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_83\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_84\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_87\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_85\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_86\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_81\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_82\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_77\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_78\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_79\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_80\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_76\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_73\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_74\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_75\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_14\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_17\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_15\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_16\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_47\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_48\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_18\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_19\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_20\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_28\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_29\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_30\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_31\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_32\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_26\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_27\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_11\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_6\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_10\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_7\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_8\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_9\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_62\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_63\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_72\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_60\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_61\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_12\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_13\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_64\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_49\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_50\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_51\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_54\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_52\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_53\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_43\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_44\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_45\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_46\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_33\ : std_logic;
signal \GNDG0\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_2\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_5\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_0\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_1\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_3\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_4\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_65\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_66\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_71\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_69\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_70\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_67\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_68\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_55\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_56\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_57\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_58\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_59\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_36\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_37\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_38\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_42\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_39\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_40\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_41\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_34\ : std_logic;
signal \generator_inst1.REGSTATZ0Z_35\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \CLK_c_g\ : std_logic;
signal \generator_inst1.REGDYN7_g\ : std_logic;
signal \RST_N_c_i_g\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \RST_N_wire\ : std_logic;
signal \SELDYN_wire\ : std_logic;
signal signal_out_wire : std_logic;
signal \SELSTAT_wire\ : std_logic;

begin
    \CLK_wire\ <= CLK;
    \RST_N_wire\ <= RST_N;
    \SELDYN_wire\ <= SELDYN;
    signal_out <= signal_out_wire;
    \SELSTAT_wire\ <= SELSTAT;

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__2334\,
            GLOBALBUFFEROUTPUT => \CLK_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2336\,
            DIN => \N__2335\,
            DOUT => \N__2334\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2336\,
            PADOUT => \N__2335\,
            PADIN => \N__2334\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RST_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2325\,
            DIN => \N__2324\,
            DOUT => \N__2323\,
            PACKAGEPIN => \RST_N_wire\
        );

    \RST_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2325\,
            PADOUT => \N__2324\,
            PADIN => \N__2323\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RST_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SELDYN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2316\,
            DIN => \N__2315\,
            DOUT => \N__2314\,
            PACKAGEPIN => \SELDYN_wire\
        );

    \SELDYN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2316\,
            PADOUT => \N__2315\,
            PADIN => \N__2314\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SELDYN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \signal_out_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2307\,
            DIN => \N__2306\,
            DOUT => \N__2305\,
            PACKAGEPIN => signal_out_wire
        );

    \signal_out_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2307\,
            PADOUT => \N__2306\,
            PADIN => \N__2305\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1418\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SELSTAT_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2298\,
            DIN => \N__2297\,
            DOUT => \N__2296\,
            PACKAGEPIN => \SELSTAT_wire\
        );

    \SELSTAT_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2298\,
            PADOUT => \N__2297\,
            PADIN => \N__2296\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SELSTAT_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__421\ : InMux
    port map (
            O => \N__2279\,
            I => \N__2276\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__2276\,
            I => \generator_inst1.REGSTATZ0Z_57\
        );

    \I__419\ : InMux
    port map (
            O => \N__2273\,
            I => \N__2270\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__2270\,
            I => \generator_inst1.REGSTATZ0Z_58\
        );

    \I__417\ : InMux
    port map (
            O => \N__2267\,
            I => \N__2264\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__2264\,
            I => \generator_inst1.REGSTATZ0Z_59\
        );

    \I__415\ : InMux
    port map (
            O => \N__2261\,
            I => \N__2258\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__2258\,
            I => \generator_inst1.REGSTATZ0Z_36\
        );

    \I__413\ : InMux
    port map (
            O => \N__2255\,
            I => \N__2252\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__2252\,
            I => \generator_inst1.REGSTATZ0Z_37\
        );

    \I__411\ : InMux
    port map (
            O => \N__2249\,
            I => \N__2246\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__2246\,
            I => \generator_inst1.REGSTATZ0Z_38\
        );

    \I__409\ : InMux
    port map (
            O => \N__2243\,
            I => \N__2240\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2240\,
            I => \generator_inst1.REGSTATZ0Z_42\
        );

    \I__407\ : InMux
    port map (
            O => \N__2237\,
            I => \N__2234\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2234\,
            I => \generator_inst1.REGSTATZ0Z_39\
        );

    \I__405\ : InMux
    port map (
            O => \N__2231\,
            I => \N__2228\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__2228\,
            I => \generator_inst1.REGSTATZ0Z_40\
        );

    \I__403\ : InMux
    port map (
            O => \N__2225\,
            I => \N__2222\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2222\,
            I => \generator_inst1.REGSTATZ0Z_41\
        );

    \I__401\ : InMux
    port map (
            O => \N__2219\,
            I => \N__2216\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__2216\,
            I => \generator_inst1.REGSTATZ0Z_34\
        );

    \I__399\ : InMux
    port map (
            O => \N__2213\,
            I => \N__2210\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__2210\,
            I => \generator_inst1.REGSTATZ0Z_35\
        );

    \I__397\ : ClkMux
    port map (
            O => \N__2207\,
            I => \N__2156\
        );

    \I__396\ : ClkMux
    port map (
            O => \N__2206\,
            I => \N__2156\
        );

    \I__395\ : ClkMux
    port map (
            O => \N__2205\,
            I => \N__2156\
        );

    \I__394\ : ClkMux
    port map (
            O => \N__2204\,
            I => \N__2156\
        );

    \I__393\ : ClkMux
    port map (
            O => \N__2203\,
            I => \N__2156\
        );

    \I__392\ : ClkMux
    port map (
            O => \N__2202\,
            I => \N__2156\
        );

    \I__391\ : ClkMux
    port map (
            O => \N__2201\,
            I => \N__2156\
        );

    \I__390\ : ClkMux
    port map (
            O => \N__2200\,
            I => \N__2156\
        );

    \I__389\ : ClkMux
    port map (
            O => \N__2199\,
            I => \N__2156\
        );

    \I__388\ : ClkMux
    port map (
            O => \N__2198\,
            I => \N__2156\
        );

    \I__387\ : ClkMux
    port map (
            O => \N__2197\,
            I => \N__2156\
        );

    \I__386\ : ClkMux
    port map (
            O => \N__2196\,
            I => \N__2156\
        );

    \I__385\ : ClkMux
    port map (
            O => \N__2195\,
            I => \N__2156\
        );

    \I__384\ : ClkMux
    port map (
            O => \N__2194\,
            I => \N__2156\
        );

    \I__383\ : ClkMux
    port map (
            O => \N__2193\,
            I => \N__2156\
        );

    \I__382\ : ClkMux
    port map (
            O => \N__2192\,
            I => \N__2156\
        );

    \I__381\ : ClkMux
    port map (
            O => \N__2191\,
            I => \N__2156\
        );

    \I__380\ : GlobalMux
    port map (
            O => \N__2156\,
            I => \N__2153\
        );

    \I__379\ : gio2CtrlBuf
    port map (
            O => \N__2153\,
            I => \CLK_c_g\
        );

    \I__378\ : CEMux
    port map (
            O => \N__2150\,
            I => \N__2108\
        );

    \I__377\ : CEMux
    port map (
            O => \N__2149\,
            I => \N__2108\
        );

    \I__376\ : CEMux
    port map (
            O => \N__2148\,
            I => \N__2108\
        );

    \I__375\ : CEMux
    port map (
            O => \N__2147\,
            I => \N__2108\
        );

    \I__374\ : CEMux
    port map (
            O => \N__2146\,
            I => \N__2108\
        );

    \I__373\ : CEMux
    port map (
            O => \N__2145\,
            I => \N__2108\
        );

    \I__372\ : CEMux
    port map (
            O => \N__2144\,
            I => \N__2108\
        );

    \I__371\ : CEMux
    port map (
            O => \N__2143\,
            I => \N__2108\
        );

    \I__370\ : CEMux
    port map (
            O => \N__2142\,
            I => \N__2108\
        );

    \I__369\ : CEMux
    port map (
            O => \N__2141\,
            I => \N__2108\
        );

    \I__368\ : CEMux
    port map (
            O => \N__2140\,
            I => \N__2108\
        );

    \I__367\ : CEMux
    port map (
            O => \N__2139\,
            I => \N__2108\
        );

    \I__366\ : CEMux
    port map (
            O => \N__2138\,
            I => \N__2108\
        );

    \I__365\ : CEMux
    port map (
            O => \N__2137\,
            I => \N__2108\
        );

    \I__364\ : GlobalMux
    port map (
            O => \N__2108\,
            I => \N__2105\
        );

    \I__363\ : gio2CtrlBuf
    port map (
            O => \N__2105\,
            I => \generator_inst1.REGDYN7_g\
        );

    \I__362\ : SRMux
    port map (
            O => \N__2102\,
            I => \N__2051\
        );

    \I__361\ : SRMux
    port map (
            O => \N__2101\,
            I => \N__2051\
        );

    \I__360\ : SRMux
    port map (
            O => \N__2100\,
            I => \N__2051\
        );

    \I__359\ : SRMux
    port map (
            O => \N__2099\,
            I => \N__2051\
        );

    \I__358\ : SRMux
    port map (
            O => \N__2098\,
            I => \N__2051\
        );

    \I__357\ : SRMux
    port map (
            O => \N__2097\,
            I => \N__2051\
        );

    \I__356\ : SRMux
    port map (
            O => \N__2096\,
            I => \N__2051\
        );

    \I__355\ : SRMux
    port map (
            O => \N__2095\,
            I => \N__2051\
        );

    \I__354\ : SRMux
    port map (
            O => \N__2094\,
            I => \N__2051\
        );

    \I__353\ : SRMux
    port map (
            O => \N__2093\,
            I => \N__2051\
        );

    \I__352\ : SRMux
    port map (
            O => \N__2092\,
            I => \N__2051\
        );

    \I__351\ : SRMux
    port map (
            O => \N__2091\,
            I => \N__2051\
        );

    \I__350\ : SRMux
    port map (
            O => \N__2090\,
            I => \N__2051\
        );

    \I__349\ : SRMux
    port map (
            O => \N__2089\,
            I => \N__2051\
        );

    \I__348\ : SRMux
    port map (
            O => \N__2088\,
            I => \N__2051\
        );

    \I__347\ : SRMux
    port map (
            O => \N__2087\,
            I => \N__2051\
        );

    \I__346\ : SRMux
    port map (
            O => \N__2086\,
            I => \N__2051\
        );

    \I__345\ : GlobalMux
    port map (
            O => \N__2051\,
            I => \N__2048\
        );

    \I__344\ : gio2CtrlBuf
    port map (
            O => \N__2048\,
            I => \RST_N_c_i_g\
        );

    \I__343\ : InMux
    port map (
            O => \N__2045\,
            I => \N__2042\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2042\,
            I => \generator_inst1.REGSTATZ0Z_66\
        );

    \I__341\ : InMux
    port map (
            O => \N__2039\,
            I => \N__2036\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2036\,
            I => \generator_inst1.REGSTATZ0Z_71\
        );

    \I__339\ : InMux
    port map (
            O => \N__2033\,
            I => \N__2030\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2030\,
            I => \generator_inst1.REGSTATZ0Z_69\
        );

    \I__337\ : InMux
    port map (
            O => \N__2027\,
            I => \N__2024\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2024\,
            I => \generator_inst1.REGSTATZ0Z_70\
        );

    \I__335\ : InMux
    port map (
            O => \N__2021\,
            I => \N__2018\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2018\,
            I => \generator_inst1.REGSTATZ0Z_67\
        );

    \I__333\ : InMux
    port map (
            O => \N__2015\,
            I => \N__2012\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2012\,
            I => \generator_inst1.REGSTATZ0Z_68\
        );

    \I__331\ : InMux
    port map (
            O => \N__2009\,
            I => \N__2006\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2006\,
            I => \generator_inst1.REGSTATZ0Z_55\
        );

    \I__329\ : InMux
    port map (
            O => \N__2003\,
            I => \N__2000\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2000\,
            I => \generator_inst1.REGSTATZ0Z_56\
        );

    \I__327\ : InMux
    port map (
            O => \N__1997\,
            I => \N__1994\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__1994\,
            I => \generator_inst1.REGSTATZ0Z_45\
        );

    \I__325\ : InMux
    port map (
            O => \N__1991\,
            I => \N__1988\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__1988\,
            I => \generator_inst1.REGSTATZ0Z_46\
        );

    \I__323\ : InMux
    port map (
            O => \N__1985\,
            I => \N__1982\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__1982\,
            I => \generator_inst1.REGSTATZ0Z_33\
        );

    \I__321\ : InMux
    port map (
            O => \N__1979\,
            I => \N__1976\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__1976\,
            I => \generator_inst1.REGSTATZ0Z_2\
        );

    \I__319\ : InMux
    port map (
            O => \N__1973\,
            I => \N__1970\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__1970\,
            I => \generator_inst1.REGSTATZ0Z_5\
        );

    \I__317\ : InMux
    port map (
            O => \N__1967\,
            I => \N__1964\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__1964\,
            I => \generator_inst1.REGSTATZ0Z_0\
        );

    \I__315\ : InMux
    port map (
            O => \N__1961\,
            I => \N__1958\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__1958\,
            I => \generator_inst1.REGSTATZ0Z_1\
        );

    \I__313\ : InMux
    port map (
            O => \N__1955\,
            I => \N__1952\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__1952\,
            I => \generator_inst1.REGSTATZ0Z_3\
        );

    \I__311\ : InMux
    port map (
            O => \N__1949\,
            I => \N__1946\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__1946\,
            I => \generator_inst1.REGSTATZ0Z_4\
        );

    \I__309\ : InMux
    port map (
            O => \N__1943\,
            I => \N__1940\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__1940\,
            I => \generator_inst1.REGSTATZ0Z_65\
        );

    \I__307\ : InMux
    port map (
            O => \N__1937\,
            I => \N__1934\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__1934\,
            I => \generator_inst1.REGSTATZ0Z_49\
        );

    \I__305\ : InMux
    port map (
            O => \N__1931\,
            I => \N__1928\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__1928\,
            I => \generator_inst1.REGSTATZ0Z_50\
        );

    \I__303\ : InMux
    port map (
            O => \N__1925\,
            I => \N__1922\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__1922\,
            I => \generator_inst1.REGSTATZ0Z_51\
        );

    \I__301\ : InMux
    port map (
            O => \N__1919\,
            I => \N__1916\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__1916\,
            I => \generator_inst1.REGSTATZ0Z_54\
        );

    \I__299\ : InMux
    port map (
            O => \N__1913\,
            I => \N__1910\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__1910\,
            I => \generator_inst1.REGSTATZ0Z_52\
        );

    \I__297\ : InMux
    port map (
            O => \N__1907\,
            I => \N__1904\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__1904\,
            I => \generator_inst1.REGSTATZ0Z_53\
        );

    \I__295\ : InMux
    port map (
            O => \N__1901\,
            I => \N__1898\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__1898\,
            I => \generator_inst1.REGSTATZ0Z_43\
        );

    \I__293\ : InMux
    port map (
            O => \N__1895\,
            I => \N__1892\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__1892\,
            I => \generator_inst1.REGSTATZ0Z_44\
        );

    \I__291\ : InMux
    port map (
            O => \N__1889\,
            I => \N__1886\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__1886\,
            I => \generator_inst1.REGSTATZ0Z_8\
        );

    \I__289\ : InMux
    port map (
            O => \N__1883\,
            I => \N__1880\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__1880\,
            I => \generator_inst1.REGSTATZ0Z_9\
        );

    \I__287\ : InMux
    port map (
            O => \N__1877\,
            I => \N__1874\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__1874\,
            I => \generator_inst1.REGSTATZ0Z_62\
        );

    \I__285\ : InMux
    port map (
            O => \N__1871\,
            I => \N__1868\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__1868\,
            I => \generator_inst1.REGSTATZ0Z_63\
        );

    \I__283\ : InMux
    port map (
            O => \N__1865\,
            I => \N__1862\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__1862\,
            I => \generator_inst1.REGSTATZ0Z_72\
        );

    \I__281\ : InMux
    port map (
            O => \N__1859\,
            I => \N__1856\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__1856\,
            I => \generator_inst1.REGSTATZ0Z_60\
        );

    \I__279\ : InMux
    port map (
            O => \N__1853\,
            I => \N__1850\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__1850\,
            I => \generator_inst1.REGSTATZ0Z_61\
        );

    \I__277\ : CascadeMux
    port map (
            O => \N__1847\,
            I => \N__1844\
        );

    \I__276\ : InMux
    port map (
            O => \N__1844\,
            I => \N__1841\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__1841\,
            I => \generator_inst1.REGSTATZ0Z_12\
        );

    \I__274\ : InMux
    port map (
            O => \N__1838\,
            I => \N__1835\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__1835\,
            I => \generator_inst1.REGSTATZ0Z_13\
        );

    \I__272\ : InMux
    port map (
            O => \N__1832\,
            I => \N__1829\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__1829\,
            I => \generator_inst1.REGSTATZ0Z_64\
        );

    \I__270\ : InMux
    port map (
            O => \N__1826\,
            I => \N__1823\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__1823\,
            I => \generator_inst1.REGSTATZ0Z_30\
        );

    \I__268\ : InMux
    port map (
            O => \N__1820\,
            I => \N__1817\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__1817\,
            I => \generator_inst1.REGSTATZ0Z_31\
        );

    \I__266\ : InMux
    port map (
            O => \N__1814\,
            I => \N__1811\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__1811\,
            I => \generator_inst1.REGSTATZ0Z_32\
        );

    \I__264\ : InMux
    port map (
            O => \N__1808\,
            I => \N__1805\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__1805\,
            I => \generator_inst1.REGSTATZ0Z_26\
        );

    \I__262\ : InMux
    port map (
            O => \N__1802\,
            I => \N__1799\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__1799\,
            I => \generator_inst1.REGSTATZ0Z_27\
        );

    \I__260\ : InMux
    port map (
            O => \N__1796\,
            I => \N__1793\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__1793\,
            I => \generator_inst1.REGSTATZ0Z_11\
        );

    \I__258\ : InMux
    port map (
            O => \N__1790\,
            I => \N__1787\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__1787\,
            I => \generator_inst1.REGSTATZ0Z_6\
        );

    \I__256\ : InMux
    port map (
            O => \N__1784\,
            I => \N__1781\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__1781\,
            I => \generator_inst1.REGSTATZ0Z_10\
        );

    \I__254\ : InMux
    port map (
            O => \N__1778\,
            I => \N__1775\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__1775\,
            I => \generator_inst1.REGSTATZ0Z_7\
        );

    \I__252\ : CascadeMux
    port map (
            O => \N__1772\,
            I => \N__1769\
        );

    \I__251\ : InMux
    port map (
            O => \N__1769\,
            I => \N__1766\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__1766\,
            I => \generator_inst1.REGSTATZ0Z_15\
        );

    \I__249\ : InMux
    port map (
            O => \N__1763\,
            I => \N__1760\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__1760\,
            I => \generator_inst1.REGSTATZ0Z_16\
        );

    \I__247\ : InMux
    port map (
            O => \N__1757\,
            I => \N__1754\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__1754\,
            I => \generator_inst1.REGSTATZ0Z_47\
        );

    \I__245\ : InMux
    port map (
            O => \N__1751\,
            I => \N__1748\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__1748\,
            I => \generator_inst1.REGSTATZ0Z_48\
        );

    \I__243\ : InMux
    port map (
            O => \N__1745\,
            I => \N__1742\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__1742\,
            I => \generator_inst1.REGSTATZ0Z_18\
        );

    \I__241\ : InMux
    port map (
            O => \N__1739\,
            I => \N__1736\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__1736\,
            I => \generator_inst1.REGSTATZ0Z_19\
        );

    \I__239\ : InMux
    port map (
            O => \N__1733\,
            I => \N__1730\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__1730\,
            I => \generator_inst1.REGSTATZ0Z_20\
        );

    \I__237\ : InMux
    port map (
            O => \N__1727\,
            I => \N__1724\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__1724\,
            I => \generator_inst1.REGSTATZ0Z_28\
        );

    \I__235\ : InMux
    port map (
            O => \N__1721\,
            I => \N__1718\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__1718\,
            I => \generator_inst1.REGSTATZ0Z_29\
        );

    \I__233\ : InMux
    port map (
            O => \N__1715\,
            I => \N__1712\
        );

    \I__232\ : LocalMux
    port map (
            O => \N__1712\,
            I => \generator_inst1.REGSTATZ0Z_79\
        );

    \I__231\ : InMux
    port map (
            O => \N__1709\,
            I => \N__1706\
        );

    \I__230\ : LocalMux
    port map (
            O => \N__1706\,
            I => \generator_inst1.REGSTATZ0Z_80\
        );

    \I__229\ : InMux
    port map (
            O => \N__1703\,
            I => \N__1700\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__1700\,
            I => \generator_inst1.REGSTATZ0Z_76\
        );

    \I__227\ : InMux
    port map (
            O => \N__1697\,
            I => \N__1694\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__1694\,
            I => \generator_inst1.REGSTATZ0Z_73\
        );

    \I__225\ : InMux
    port map (
            O => \N__1691\,
            I => \N__1688\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__1688\,
            I => \generator_inst1.REGSTATZ0Z_74\
        );

    \I__223\ : InMux
    port map (
            O => \N__1685\,
            I => \N__1682\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__1682\,
            I => \generator_inst1.REGSTATZ0Z_75\
        );

    \I__221\ : InMux
    port map (
            O => \N__1679\,
            I => \N__1676\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__1676\,
            I => \generator_inst1.REGSTATZ0Z_14\
        );

    \I__219\ : InMux
    port map (
            O => \N__1673\,
            I => \N__1670\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__1670\,
            I => \generator_inst1.REGSTATZ0Z_17\
        );

    \I__217\ : InMux
    port map (
            O => \N__1667\,
            I => \N__1664\
        );

    \I__216\ : LocalMux
    port map (
            O => \N__1664\,
            I => \generator_inst1.REGSTATZ0Z_83\
        );

    \I__215\ : InMux
    port map (
            O => \N__1661\,
            I => \N__1658\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__1658\,
            I => \generator_inst1.REGSTATZ0Z_84\
        );

    \I__213\ : InMux
    port map (
            O => \N__1655\,
            I => \N__1652\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__1652\,
            I => \generator_inst1.REGSTATZ0Z_87\
        );

    \I__211\ : InMux
    port map (
            O => \N__1649\,
            I => \N__1646\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__1646\,
            I => \generator_inst1.REGSTATZ0Z_85\
        );

    \I__209\ : InMux
    port map (
            O => \N__1643\,
            I => \N__1640\
        );

    \I__208\ : LocalMux
    port map (
            O => \N__1640\,
            I => \generator_inst1.REGSTATZ0Z_86\
        );

    \I__207\ : InMux
    port map (
            O => \N__1637\,
            I => \N__1634\
        );

    \I__206\ : LocalMux
    port map (
            O => \N__1634\,
            I => \generator_inst1.REGSTATZ0Z_81\
        );

    \I__205\ : InMux
    port map (
            O => \N__1631\,
            I => \N__1628\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__1628\,
            I => \generator_inst1.REGSTATZ0Z_82\
        );

    \I__203\ : InMux
    port map (
            O => \N__1625\,
            I => \N__1622\
        );

    \I__202\ : LocalMux
    port map (
            O => \N__1622\,
            I => \generator_inst1.REGSTATZ0Z_77\
        );

    \I__201\ : InMux
    port map (
            O => \N__1619\,
            I => \N__1616\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__1616\,
            I => \generator_inst1.REGSTATZ0Z_78\
        );

    \I__199\ : InMux
    port map (
            O => \N__1613\,
            I => \N__1610\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__1610\,
            I => \generator_inst1.REGDYNZ0Z_0\
        );

    \I__197\ : InMux
    port map (
            O => \N__1607\,
            I => \N__1604\
        );

    \I__196\ : LocalMux
    port map (
            O => \N__1604\,
            I => \generator_inst1.REGSTATZ0Z_24\
        );

    \I__195\ : InMux
    port map (
            O => \N__1601\,
            I => \N__1598\
        );

    \I__194\ : LocalMux
    port map (
            O => \N__1598\,
            I => \generator_inst1.REGSTATZ0Z_25\
        );

    \I__193\ : InMux
    port map (
            O => \N__1595\,
            I => \N__1592\
        );

    \I__192\ : LocalMux
    port map (
            O => \N__1592\,
            I => \generator_inst1.REGSTATZ0Z_22\
        );

    \I__191\ : InMux
    port map (
            O => \N__1589\,
            I => \N__1586\
        );

    \I__190\ : LocalMux
    port map (
            O => \N__1586\,
            I => \generator_inst1.REGSTATZ0Z_23\
        );

    \I__189\ : InMux
    port map (
            O => \N__1583\,
            I => \N__1580\
        );

    \I__188\ : LocalMux
    port map (
            O => \N__1580\,
            I => \generator_inst1.REGSTATZ0Z_21\
        );

    \I__187\ : InMux
    port map (
            O => \N__1577\,
            I => \N__1574\
        );

    \I__186\ : LocalMux
    port map (
            O => \N__1574\,
            I => \N__1571\
        );

    \I__185\ : IoSpan4Mux
    port map (
            O => \N__1571\,
            I => \N__1567\
        );

    \I__184\ : InMux
    port map (
            O => \N__1570\,
            I => \N__1564\
        );

    \I__183\ : Odrv4
    port map (
            O => \N__1567\,
            I => \SELSTAT_c\
        );

    \I__182\ : LocalMux
    port map (
            O => \N__1564\,
            I => \SELSTAT_c\
        );

    \I__181\ : InMux
    port map (
            O => \N__1559\,
            I => \N__1556\
        );

    \I__180\ : LocalMux
    port map (
            O => \N__1556\,
            I => \N__1552\
        );

    \I__179\ : CEMux
    port map (
            O => \N__1555\,
            I => \N__1549\
        );

    \I__178\ : Span4Mux_h
    port map (
            O => \N__1552\,
            I => \N__1544\
        );

    \I__177\ : LocalMux
    port map (
            O => \N__1549\,
            I => \N__1544\
        );

    \I__176\ : Span4Mux_v
    port map (
            O => \N__1544\,
            I => \N__1540\
        );

    \I__175\ : CEMux
    port map (
            O => \N__1543\,
            I => \N__1537\
        );

    \I__174\ : Span4Mux_v
    port map (
            O => \N__1540\,
            I => \N__1531\
        );

    \I__173\ : LocalMux
    port map (
            O => \N__1537\,
            I => \N__1531\
        );

    \I__172\ : InMux
    port map (
            O => \N__1536\,
            I => \N__1528\
        );

    \I__171\ : Span4Mux_v
    port map (
            O => \N__1531\,
            I => \N__1523\
        );

    \I__170\ : LocalMux
    port map (
            O => \N__1528\,
            I => \N__1523\
        );

    \I__169\ : Span4Mux_v
    port map (
            O => \N__1523\,
            I => \N__1520\
        );

    \I__168\ : Odrv4
    port map (
            O => \N__1520\,
            I => \SELDYN_c\
        );

    \I__167\ : IoInMux
    port map (
            O => \N__1517\,
            I => \N__1514\
        );

    \I__166\ : LocalMux
    port map (
            O => \N__1514\,
            I => \generator_inst1.REGDYNZ0Z7\
        );

    \I__165\ : InMux
    port map (
            O => \N__1511\,
            I => \N__1508\
        );

    \I__164\ : LocalMux
    port map (
            O => \N__1508\,
            I => \generator_inst1.REGDYNZ0Z_11\
        );

    \I__163\ : InMux
    port map (
            O => \N__1505\,
            I => \N__1502\
        );

    \I__162\ : LocalMux
    port map (
            O => \N__1502\,
            I => \generator_inst1.REGDYNZ0Z_9\
        );

    \I__161\ : InMux
    port map (
            O => \N__1499\,
            I => \N__1496\
        );

    \I__160\ : LocalMux
    port map (
            O => \N__1496\,
            I => \generator_inst1.REGDYNZ0Z_10\
        );

    \I__159\ : InMux
    port map (
            O => \N__1493\,
            I => \N__1490\
        );

    \I__158\ : LocalMux
    port map (
            O => \N__1490\,
            I => \generator_inst1.REGDYNZ0Z_1\
        );

    \I__157\ : InMux
    port map (
            O => \N__1487\,
            I => \N__1484\
        );

    \I__156\ : LocalMux
    port map (
            O => \N__1484\,
            I => \generator_inst1.REGDYNZ0Z_2\
        );

    \I__155\ : InMux
    port map (
            O => \N__1481\,
            I => \N__1478\
        );

    \I__154\ : LocalMux
    port map (
            O => \N__1478\,
            I => \generator_inst1.REGDYNZ0Z_6\
        );

    \I__153\ : InMux
    port map (
            O => \N__1475\,
            I => \N__1472\
        );

    \I__152\ : LocalMux
    port map (
            O => \N__1472\,
            I => \generator_inst1.REGDYNZ0Z_7\
        );

    \I__151\ : InMux
    port map (
            O => \N__1469\,
            I => \N__1466\
        );

    \I__150\ : LocalMux
    port map (
            O => \N__1466\,
            I => \generator_inst1.REGDYNZ0Z_5\
        );

    \I__149\ : InMux
    port map (
            O => \N__1463\,
            I => \N__1460\
        );

    \I__148\ : LocalMux
    port map (
            O => \N__1460\,
            I => \generator_inst1.REGDYNZ0Z_3\
        );

    \I__147\ : InMux
    port map (
            O => \N__1457\,
            I => \N__1454\
        );

    \I__146\ : LocalMux
    port map (
            O => \N__1454\,
            I => \generator_inst1.REGDYNZ0Z_4\
        );

    \I__145\ : InMux
    port map (
            O => \N__1451\,
            I => \N__1448\
        );

    \I__144\ : LocalMux
    port map (
            O => \N__1448\,
            I => \N__1445\
        );

    \I__143\ : Span4Mux_v
    port map (
            O => \N__1445\,
            I => \N__1442\
        );

    \I__142\ : Odrv4
    port map (
            O => \N__1442\,
            I => \RST_N_c\
        );

    \I__141\ : IoInMux
    port map (
            O => \N__1439\,
            I => \N__1436\
        );

    \I__140\ : LocalMux
    port map (
            O => \N__1436\,
            I => \N__1433\
        );

    \I__139\ : Span4Mux_s0_h
    port map (
            O => \N__1433\,
            I => \N__1430\
        );

    \I__138\ : Span4Mux_v
    port map (
            O => \N__1430\,
            I => \N__1427\
        );

    \I__137\ : Odrv4
    port map (
            O => \N__1427\,
            I => \RST_N_c_i\
        );

    \I__136\ : InMux
    port map (
            O => \N__1424\,
            I => \N__1421\
        );

    \I__135\ : LocalMux
    port map (
            O => \N__1421\,
            I => generated_signal
        );

    \I__134\ : IoInMux
    port map (
            O => \N__1418\,
            I => \N__1415\
        );

    \I__133\ : LocalMux
    port map (
            O => \N__1415\,
            I => \N__1412\
        );

    \I__132\ : IoSpan4Mux
    port map (
            O => \N__1412\,
            I => \N__1409\
        );

    \I__131\ : IoSpan4Mux
    port map (
            O => \N__1409\,
            I => \N__1406\
        );

    \I__130\ : IoSpan4Mux
    port map (
            O => \N__1406\,
            I => \N__1403\
        );

    \I__129\ : Odrv4
    port map (
            O => \N__1403\,
            I => signal_out_c
        );

    \I__128\ : InMux
    port map (
            O => \N__1400\,
            I => \N__1397\
        );

    \I__127\ : LocalMux
    port map (
            O => \N__1397\,
            I => \generator_inst1.REGDYNZ0Z_8\
        );

    \I__126\ : InMux
    port map (
            O => \N__1394\,
            I => \N__1391\
        );

    \I__125\ : LocalMux
    port map (
            O => \N__1391\,
            I => \generator_inst1.REGDYNZ0Z_12\
        );

    \I__124\ : InMux
    port map (
            O => \N__1388\,
            I => \N__1385\
        );

    \I__123\ : LocalMux
    port map (
            O => \N__1385\,
            I => \generator_inst1.REGDYNZ0Z_13\
        );

    \I__122\ : InMux
    port map (
            O => \N__1382\,
            I => \N__1379\
        );

    \I__121\ : LocalMux
    port map (
            O => \N__1379\,
            I => \generator_inst1.REGDYNZ0Z_14\
        );

    \I__120\ : CascadeMux
    port map (
            O => \N__1376\,
            I => \N__1373\
        );

    \I__119\ : InMux
    port map (
            O => \N__1373\,
            I => \N__1370\
        );

    \I__118\ : LocalMux
    port map (
            O => \N__1370\,
            I => \generator_inst1.REGDYNZ0Z_15\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \generator_inst1.REGDYN7_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__1517\,
            GLOBALBUFFEROUTPUT => \generator_inst1.REGDYN7_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \RST_N_ibuf_RNIBJGC_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__1439\,
            GLOBALBUFFEROUTPUT => \RST_N_c_i_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \RST_N_ibuf_RNIBJGC_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1451\,
            lcout => \RST_N_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.signal_out_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110010000100000"
        )
    port map (
            in0 => \N__1577\,
            in1 => \N__1559\,
            in2 => \N__1376\,
            in3 => \N__1655\,
            lcout => generated_signal,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2200\,
            ce => 'H',
            sr => \N__2095\
        );

    \receptor_inst1.signal_out_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1424\,
            lcout => signal_out_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2200\,
            ce => 'H',
            sr => \N__2095\
        );

    \generator_inst1.REGDYN_9_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1400\,
            lcout => \generator_inst1.REGDYNZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2196\,
            ce => \N__1555\,
            sr => \N__2092\
        );

    \generator_inst1.REGDYN_8_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1475\,
            lcout => \generator_inst1.REGDYNZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2196\,
            ce => \N__1555\,
            sr => \N__2092\
        );

    \generator_inst1.REGDYN_12_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1511\,
            lcout => \generator_inst1.REGDYNZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2196\,
            ce => \N__1555\,
            sr => \N__2092\
        );

    \generator_inst1.REGDYN_13_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1394\,
            lcout => \generator_inst1.REGDYNZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2196\,
            ce => \N__1555\,
            sr => \N__2092\
        );

    \generator_inst1.REGDYN_14_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1388\,
            lcout => \generator_inst1.REGDYNZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2196\,
            ce => \N__1555\,
            sr => \N__2092\
        );

    \generator_inst1.REGDYN_15_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1382\,
            lcout => \generator_inst1.REGDYNZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2196\,
            ce => \N__1555\,
            sr => \N__2092\
        );

    \generator_inst1.REGDYN_11_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1499\,
            lcout => \generator_inst1.REGDYNZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2196\,
            ce => \N__1555\,
            sr => \N__2092\
        );

    \generator_inst1.REGDYN_10_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1505\,
            lcout => \generator_inst1.REGDYNZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2196\,
            ce => \N__1555\,
            sr => \N__2092\
        );

    \generator_inst1.REGDYN_1_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1613\,
            lcout => \generator_inst1.REGDYNZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2193\,
            ce => \N__1543\,
            sr => \N__2089\
        );

    \generator_inst1.REGDYN_2_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1493\,
            lcout => \generator_inst1.REGDYNZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2193\,
            ce => \N__1543\,
            sr => \N__2089\
        );

    \generator_inst1.REGDYN_3_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1487\,
            lcout => \generator_inst1.REGDYNZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2193\,
            ce => \N__1543\,
            sr => \N__2089\
        );

    \generator_inst1.REGDYN_6_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1469\,
            lcout => \generator_inst1.REGDYNZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2193\,
            ce => \N__1543\,
            sr => \N__2089\
        );

    \generator_inst1.REGDYN_7_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1481\,
            lcout => \generator_inst1.REGDYNZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2193\,
            ce => \N__1543\,
            sr => \N__2089\
        );

    \generator_inst1.REGDYN_5_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1457\,
            lcout => \generator_inst1.REGDYNZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2193\,
            ce => \N__1543\,
            sr => \N__2089\
        );

    \generator_inst1.REGDYN_4_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1463\,
            lcout => \generator_inst1.REGDYNZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2193\,
            ce => \N__1543\,
            sr => \N__2089\
        );

    \generator_inst1.REGDYN_0_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \generator_inst1.REGDYNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2193\,
            ce => \N__1543\,
            sr => \N__2089\
        );

    \generator_inst1.REGSTAT_24_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1589\,
            lcout => \generator_inst1.REGSTATZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2191\,
            ce => \N__2137\,
            sr => \N__2087\
        );

    \generator_inst1.REGSTAT_26_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1601\,
            lcout => \generator_inst1.REGSTATZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2191\,
            ce => \N__2137\,
            sr => \N__2087\
        );

    \generator_inst1.REGSTAT_25_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1607\,
            lcout => \generator_inst1.REGSTATZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2191\,
            ce => \N__2137\,
            sr => \N__2087\
        );

    \generator_inst1.REGSTAT_22_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1583\,
            lcout => \generator_inst1.REGSTATZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2191\,
            ce => \N__2137\,
            sr => \N__2087\
        );

    \generator_inst1.REGSTAT_23_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1595\,
            lcout => \generator_inst1.REGSTATZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2191\,
            ce => \N__2137\,
            sr => \N__2087\
        );

    \generator_inst1.REGSTAT_21_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1733\,
            lcout => \generator_inst1.REGSTATZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2191\,
            ce => \N__2137\,
            sr => \N__2087\
        );

    \generator_inst1.REGDYN7_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__1570\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1536\,
            lcout => \generator_inst1.REGDYNZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.REGSTAT_83_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1631\,
            lcout => \generator_inst1.REGSTATZ0Z_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2204\,
            ce => \N__2147\,
            sr => \N__2099\
        );

    \generator_inst1.REGSTAT_84_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1667\,
            lcout => \generator_inst1.REGSTATZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2204\,
            ce => \N__2147\,
            sr => \N__2099\
        );

    \generator_inst1.REGSTAT_81_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1709\,
            lcout => \generator_inst1.REGSTATZ0Z_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2204\,
            ce => \N__2147\,
            sr => \N__2099\
        );

    \generator_inst1.REGSTAT_85_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1661\,
            lcout => \generator_inst1.REGSTATZ0Z_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2204\,
            ce => \N__2147\,
            sr => \N__2099\
        );

    \generator_inst1.REGSTAT_87_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1643\,
            lcout => \generator_inst1.REGSTATZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2204\,
            ce => \N__2147\,
            sr => \N__2099\
        );

    \generator_inst1.REGSTAT_86_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1649\,
            lcout => \generator_inst1.REGSTATZ0Z_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2204\,
            ce => \N__2147\,
            sr => \N__2099\
        );

    \generator_inst1.REGSTAT_82_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1637\,
            lcout => \generator_inst1.REGSTATZ0Z_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2204\,
            ce => \N__2147\,
            sr => \N__2099\
        );

    \generator_inst1.REGSTAT_79_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1619\,
            lcout => \generator_inst1.REGSTATZ0Z_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2201\,
            ce => \N__2144\,
            sr => \N__2096\
        );

    \generator_inst1.REGSTAT_77_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1703\,
            lcout => \generator_inst1.REGSTATZ0Z_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2201\,
            ce => \N__2144\,
            sr => \N__2096\
        );

    \generator_inst1.REGSTAT_78_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1625\,
            lcout => \generator_inst1.REGSTATZ0Z_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2201\,
            ce => \N__2144\,
            sr => \N__2096\
        );

    \generator_inst1.REGSTAT_80_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1715\,
            lcout => \generator_inst1.REGSTATZ0Z_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2201\,
            ce => \N__2144\,
            sr => \N__2096\
        );

    \generator_inst1.REGSTAT_15_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1679\,
            lcout => \generator_inst1.REGSTATZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2197\,
            ce => \N__2141\,
            sr => \N__2093\
        );

    \generator_inst1.REGSTAT_76_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1685\,
            lcout => \generator_inst1.REGSTATZ0Z_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2197\,
            ce => \N__2141\,
            sr => \N__2093\
        );

    \generator_inst1.REGSTAT_74_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1697\,
            lcout => \generator_inst1.REGSTATZ0Z_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2197\,
            ce => \N__2141\,
            sr => \N__2093\
        );

    \generator_inst1.REGSTAT_73_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1865\,
            lcout => \generator_inst1.REGSTATZ0Z_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2197\,
            ce => \N__2141\,
            sr => \N__2093\
        );

    \generator_inst1.REGSTAT_75_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1691\,
            lcout => \generator_inst1.REGSTATZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2197\,
            ce => \N__2141\,
            sr => \N__2093\
        );

    \generator_inst1.REGSTAT_14_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1838\,
            lcout => \generator_inst1.REGSTATZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2197\,
            ce => \N__2141\,
            sr => \N__2093\
        );

    \generator_inst1.REGSTAT_17_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1763\,
            lcout => \generator_inst1.REGSTATZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2194\,
            ce => \N__2139\,
            sr => \N__2090\
        );

    \generator_inst1.REGSTAT_18_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1673\,
            lcout => \generator_inst1.REGSTATZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2194\,
            ce => \N__2139\,
            sr => \N__2090\
        );

    \generator_inst1.REGSTAT_47_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1991\,
            lcout => \generator_inst1.REGSTATZ0Z_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2194\,
            ce => \N__2139\,
            sr => \N__2090\
        );

    \generator_inst1.REGSTAT_49_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1751\,
            lcout => \generator_inst1.REGSTATZ0Z_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2194\,
            ce => \N__2139\,
            sr => \N__2090\
        );

    \generator_inst1.REGSTAT_16_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1772\,
            in3 => \_gnd_net_\,
            lcout => \generator_inst1.REGSTATZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2194\,
            ce => \N__2139\,
            sr => \N__2090\
        );

    \generator_inst1.REGSTAT_48_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1757\,
            lcout => \generator_inst1.REGSTATZ0Z_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2194\,
            ce => \N__2139\,
            sr => \N__2090\
        );

    \generator_inst1.REGSTAT_19_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1745\,
            lcout => \generator_inst1.REGSTATZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2194\,
            ce => \N__2139\,
            sr => \N__2090\
        );

    \generator_inst1.REGSTAT_20_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1739\,
            lcout => \generator_inst1.REGSTATZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2194\,
            ce => \N__2139\,
            sr => \N__2090\
        );

    \generator_inst1.REGSTAT_33_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1814\,
            lcout => \generator_inst1.REGSTATZ0Z_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2192\,
            ce => \N__2138\,
            sr => \N__2086\
        );

    \generator_inst1.REGSTAT_28_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1802\,
            lcout => \generator_inst1.REGSTATZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2192\,
            ce => \N__2138\,
            sr => \N__2086\
        );

    \generator_inst1.REGSTAT_29_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1727\,
            lcout => \generator_inst1.REGSTATZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2192\,
            ce => \N__2138\,
            sr => \N__2086\
        );

    \generator_inst1.REGSTAT_30_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1721\,
            lcout => \generator_inst1.REGSTATZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2192\,
            ce => \N__2138\,
            sr => \N__2086\
        );

    \generator_inst1.REGSTAT_31_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1826\,
            lcout => \generator_inst1.REGSTATZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2192\,
            ce => \N__2138\,
            sr => \N__2086\
        );

    \generator_inst1.REGSTAT_32_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1820\,
            lcout => \generator_inst1.REGSTATZ0Z_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2192\,
            ce => \N__2138\,
            sr => \N__2086\
        );

    \generator_inst1.REGSTAT_27_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1808\,
            lcout => \generator_inst1.REGSTATZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2192\,
            ce => \N__2138\,
            sr => \N__2086\
        );

    \generator_inst1.REGSTAT_11_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1784\,
            lcout => \generator_inst1.REGSTATZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2205\,
            ce => \N__2148\,
            sr => \N__2100\
        );

    \generator_inst1.REGSTAT_12_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1796\,
            lcout => \generator_inst1.REGSTATZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2205\,
            ce => \N__2148\,
            sr => \N__2100\
        );

    \generator_inst1.REGSTAT_7_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1790\,
            lcout => \generator_inst1.REGSTATZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2205\,
            ce => \N__2148\,
            sr => \N__2100\
        );

    \generator_inst1.REGSTAT_6_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1973\,
            lcout => \generator_inst1.REGSTATZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2205\,
            ce => \N__2148\,
            sr => \N__2100\
        );

    \generator_inst1.REGSTAT_10_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1883\,
            lcout => \generator_inst1.REGSTATZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2205\,
            ce => \N__2148\,
            sr => \N__2100\
        );

    \generator_inst1.REGSTAT_8_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1778\,
            lcout => \generator_inst1.REGSTATZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2205\,
            ce => \N__2148\,
            sr => \N__2100\
        );

    \generator_inst1.REGSTAT_9_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1889\,
            lcout => \generator_inst1.REGSTATZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2205\,
            ce => \N__2148\,
            sr => \N__2100\
        );

    \generator_inst1.REGSTAT_62_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1853\,
            lcout => \generator_inst1.REGSTATZ0Z_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2202\,
            ce => \N__2145\,
            sr => \N__2097\
        );

    \generator_inst1.REGSTAT_64_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1871\,
            lcout => \generator_inst1.REGSTATZ0Z_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2202\,
            ce => \N__2145\,
            sr => \N__2097\
        );

    \generator_inst1.REGSTAT_63_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1877\,
            lcout => \generator_inst1.REGSTATZ0Z_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2202\,
            ce => \N__2145\,
            sr => \N__2097\
        );

    \generator_inst1.REGSTAT_60_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2267\,
            lcout => \generator_inst1.REGSTATZ0Z_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2202\,
            ce => \N__2145\,
            sr => \N__2097\
        );

    \generator_inst1.REGSTAT_72_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2039\,
            lcout => \generator_inst1.REGSTATZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2202\,
            ce => \N__2145\,
            sr => \N__2097\
        );

    \generator_inst1.REGSTAT_61_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1859\,
            lcout => \generator_inst1.REGSTATZ0Z_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2202\,
            ce => \N__2145\,
            sr => \N__2097\
        );

    \generator_inst1.REGSTAT_13_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1847\,
            in3 => \_gnd_net_\,
            lcout => \generator_inst1.REGSTATZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2202\,
            ce => \N__2145\,
            sr => \N__2097\
        );

    \generator_inst1.REGSTAT_65_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1832\,
            lcout => \generator_inst1.REGSTATZ0Z_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2202\,
            ce => \N__2145\,
            sr => \N__2097\
        );

    \generator_inst1.REGSTAT_55_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1919\,
            lcout => \generator_inst1.REGSTATZ0Z_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2198\,
            ce => \N__2142\,
            sr => \N__2094\
        );

    \generator_inst1.REGSTAT_50_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1937\,
            lcout => \generator_inst1.REGSTATZ0Z_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2198\,
            ce => \N__2142\,
            sr => \N__2094\
        );

    \generator_inst1.REGSTAT_51_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1931\,
            lcout => \generator_inst1.REGSTATZ0Z_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2198\,
            ce => \N__2142\,
            sr => \N__2094\
        );

    \generator_inst1.REGSTAT_52_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1925\,
            lcout => \generator_inst1.REGSTATZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2198\,
            ce => \N__2142\,
            sr => \N__2094\
        );

    \generator_inst1.REGSTAT_54_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1907\,
            lcout => \generator_inst1.REGSTATZ0Z_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2198\,
            ce => \N__2142\,
            sr => \N__2094\
        );

    \generator_inst1.REGSTAT_53_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1913\,
            lcout => \generator_inst1.REGSTATZ0Z_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2198\,
            ce => \N__2142\,
            sr => \N__2094\
        );

    \generator_inst1.REGSTAT_43_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2243\,
            lcout => \generator_inst1.REGSTATZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2195\,
            ce => \N__2140\,
            sr => \N__2088\
        );

    \generator_inst1.REGSTAT_44_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1901\,
            lcout => \generator_inst1.REGSTATZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2195\,
            ce => \N__2140\,
            sr => \N__2088\
        );

    \generator_inst1.REGSTAT_45_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1895\,
            lcout => \generator_inst1.REGSTATZ0Z_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2195\,
            ce => \N__2140\,
            sr => \N__2088\
        );

    \generator_inst1.REGSTAT_46_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1997\,
            lcout => \generator_inst1.REGSTATZ0Z_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2195\,
            ce => \N__2140\,
            sr => \N__2088\
        );

    \generator_inst1.REGSTAT_34_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1985\,
            lcout => \generator_inst1.REGSTATZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2195\,
            ce => \N__2140\,
            sr => \N__2088\
        );

    \generator_inst1.REGSTAT_0_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \generator_inst1.REGSTATZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2207\,
            ce => \N__2150\,
            sr => \N__2102\
        );

    \generator_inst1.REGSTAT_2_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1961\,
            lcout => \generator_inst1.REGSTATZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2207\,
            ce => \N__2150\,
            sr => \N__2102\
        );

    \generator_inst1.REGSTAT_3_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1979\,
            lcout => \generator_inst1.REGSTATZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2207\,
            ce => \N__2150\,
            sr => \N__2102\
        );

    \generator_inst1.REGSTAT_5_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1949\,
            lcout => \generator_inst1.REGSTATZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2207\,
            ce => \N__2150\,
            sr => \N__2102\
        );

    \generator_inst1.REGSTAT_1_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1967\,
            lcout => \generator_inst1.REGSTATZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2207\,
            ce => \N__2150\,
            sr => \N__2102\
        );

    \generator_inst1.REGSTAT_4_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1955\,
            lcout => \generator_inst1.REGSTATZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2207\,
            ce => \N__2150\,
            sr => \N__2102\
        );

    \generator_inst1.REGSTAT_66_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1943\,
            lcout => \generator_inst1.REGSTATZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2206\,
            ce => \N__2149\,
            sr => \N__2101\
        );

    \generator_inst1.REGSTAT_67_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2045\,
            lcout => \generator_inst1.REGSTATZ0Z_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2206\,
            ce => \N__2149\,
            sr => \N__2101\
        );

    \generator_inst1.REGSTAT_69_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2015\,
            lcout => \generator_inst1.REGSTATZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2206\,
            ce => \N__2149\,
            sr => \N__2101\
        );

    \generator_inst1.REGSTAT_71_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2027\,
            lcout => \generator_inst1.REGSTATZ0Z_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2206\,
            ce => \N__2149\,
            sr => \N__2101\
        );

    \generator_inst1.REGSTAT_70_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2033\,
            lcout => \generator_inst1.REGSTATZ0Z_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2206\,
            ce => \N__2149\,
            sr => \N__2101\
        );

    \generator_inst1.REGSTAT_68_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2021\,
            lcout => \generator_inst1.REGSTATZ0Z_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2206\,
            ce => \N__2149\,
            sr => \N__2101\
        );

    \generator_inst1.REGSTAT_56_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2009\,
            lcout => \generator_inst1.REGSTATZ0Z_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2203\,
            ce => \N__2146\,
            sr => \N__2098\
        );

    \generator_inst1.REGSTAT_57_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2003\,
            lcout => \generator_inst1.REGSTATZ0Z_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2203\,
            ce => \N__2146\,
            sr => \N__2098\
        );

    \generator_inst1.REGSTAT_36_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2213\,
            lcout => \generator_inst1.REGSTATZ0Z_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2203\,
            ce => \N__2146\,
            sr => \N__2098\
        );

    \generator_inst1.REGSTAT_38_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2255\,
            lcout => \generator_inst1.REGSTATZ0Z_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2203\,
            ce => \N__2146\,
            sr => \N__2098\
        );

    \generator_inst1.REGSTAT_58_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2279\,
            lcout => \generator_inst1.REGSTATZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2203\,
            ce => \N__2146\,
            sr => \N__2098\
        );

    \generator_inst1.REGSTAT_59_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2273\,
            lcout => \generator_inst1.REGSTATZ0Z_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2203\,
            ce => \N__2146\,
            sr => \N__2098\
        );

    \generator_inst1.REGSTAT_37_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2261\,
            lcout => \generator_inst1.REGSTATZ0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2203\,
            ce => \N__2146\,
            sr => \N__2098\
        );

    \generator_inst1.REGSTAT_39_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2249\,
            lcout => \generator_inst1.REGSTATZ0Z_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2199\,
            ce => \N__2143\,
            sr => \N__2091\
        );

    \generator_inst1.REGSTAT_42_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2225\,
            lcout => \generator_inst1.REGSTATZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2199\,
            ce => \N__2143\,
            sr => \N__2091\
        );

    \generator_inst1.REGSTAT_40_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2237\,
            lcout => \generator_inst1.REGSTATZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2199\,
            ce => \N__2143\,
            sr => \N__2091\
        );

    \generator_inst1.REGSTAT_41_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2231\,
            lcout => \generator_inst1.REGSTATZ0Z_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2199\,
            ce => \N__2143\,
            sr => \N__2091\
        );

    \generator_inst1.REGSTAT_35_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2219\,
            lcout => \generator_inst1.REGSTATZ0Z_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2199\,
            ce => \N__2143\,
            sr => \N__2091\
        );
end \INTERFACE\;
