-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 18 2025 09:13:17

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    generated_signal : out std_logic;
    RST_N : in std_logic;
    ENdin : out std_logic;
    CLK : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__1628\ : std_logic;
signal \N__1627\ : std_logic;
signal \N__1626\ : std_logic;
signal \N__1617\ : std_logic;
signal \N__1616\ : std_logic;
signal \N__1615\ : std_logic;
signal \N__1608\ : std_logic;
signal \N__1607\ : std_logic;
signal \N__1606\ : std_logic;
signal \N__1599\ : std_logic;
signal \N__1598\ : std_logic;
signal \N__1597\ : std_logic;
signal \N__1580\ : std_logic;
signal \N__1579\ : std_logic;
signal \N__1578\ : std_logic;
signal \N__1575\ : std_logic;
signal \N__1572\ : std_logic;
signal \N__1569\ : std_logic;
signal \N__1564\ : std_logic;
signal \N__1561\ : std_logic;
signal \N__1556\ : std_logic;
signal \N__1553\ : std_logic;
signal \N__1552\ : std_logic;
signal \N__1551\ : std_logic;
signal \N__1548\ : std_logic;
signal \N__1545\ : std_logic;
signal \N__1542\ : std_logic;
signal \N__1535\ : std_logic;
signal \N__1532\ : std_logic;
signal \N__1531\ : std_logic;
signal \N__1528\ : std_logic;
signal \N__1525\ : std_logic;
signal \N__1520\ : std_logic;
signal \N__1517\ : std_logic;
signal \N__1516\ : std_logic;
signal \N__1515\ : std_logic;
signal \N__1512\ : std_logic;
signal \N__1507\ : std_logic;
signal \N__1504\ : std_logic;
signal \N__1499\ : std_logic;
signal \N__1496\ : std_logic;
signal \N__1495\ : std_logic;
signal \N__1492\ : std_logic;
signal \N__1489\ : std_logic;
signal \N__1484\ : std_logic;
signal \N__1481\ : std_logic;
signal \N__1478\ : std_logic;
signal \N__1477\ : std_logic;
signal \N__1474\ : std_logic;
signal \N__1471\ : std_logic;
signal \N__1468\ : std_logic;
signal \N__1463\ : std_logic;
signal \N__1460\ : std_logic;
signal \N__1459\ : std_logic;
signal \N__1458\ : std_logic;
signal \N__1457\ : std_logic;
signal \N__1456\ : std_logic;
signal \N__1455\ : std_logic;
signal \N__1454\ : std_logic;
signal \N__1453\ : std_logic;
signal \N__1444\ : std_logic;
signal \N__1435\ : std_logic;
signal \N__1430\ : std_logic;
signal \N__1427\ : std_logic;
signal \N__1426\ : std_logic;
signal \N__1423\ : std_logic;
signal \N__1420\ : std_logic;
signal \N__1415\ : std_logic;
signal \N__1414\ : std_logic;
signal \N__1413\ : std_logic;
signal \N__1412\ : std_logic;
signal \N__1411\ : std_logic;
signal \N__1410\ : std_logic;
signal \N__1409\ : std_logic;
signal \N__1408\ : std_logic;
signal \N__1407\ : std_logic;
signal \N__1406\ : std_logic;
signal \N__1405\ : std_logic;
signal \N__1404\ : std_logic;
signal \N__1379\ : std_logic;
signal \N__1376\ : std_logic;
signal \N__1373\ : std_logic;
signal \N__1372\ : std_logic;
signal \N__1371\ : std_logic;
signal \N__1370\ : std_logic;
signal \N__1369\ : std_logic;
signal \N__1368\ : std_logic;
signal \N__1367\ : std_logic;
signal \N__1366\ : std_logic;
signal \N__1365\ : std_logic;
signal \N__1346\ : std_logic;
signal \N__1343\ : std_logic;
signal \N__1340\ : std_logic;
signal \N__1339\ : std_logic;
signal \N__1336\ : std_logic;
signal \N__1333\ : std_logic;
signal \N__1328\ : std_logic;
signal \N__1325\ : std_logic;
signal \N__1322\ : std_logic;
signal \N__1319\ : std_logic;
signal \N__1316\ : std_logic;
signal \N__1315\ : std_logic;
signal \N__1314\ : std_logic;
signal \N__1313\ : std_logic;
signal \N__1312\ : std_logic;
signal \N__1311\ : std_logic;
signal \N__1310\ : std_logic;
signal \N__1309\ : std_logic;
signal \N__1308\ : std_logic;
signal \N__1307\ : std_logic;
signal \N__1306\ : std_logic;
signal \N__1305\ : std_logic;
signal \N__1304\ : std_logic;
signal \N__1303\ : std_logic;
signal \N__1302\ : std_logic;
signal \N__1299\ : std_logic;
signal \N__1286\ : std_logic;
signal \N__1269\ : std_logic;
signal \N__1262\ : std_logic;
signal \N__1261\ : std_logic;
signal \N__1260\ : std_logic;
signal \N__1259\ : std_logic;
signal \N__1256\ : std_logic;
signal \N__1253\ : std_logic;
signal \N__1248\ : std_logic;
signal \N__1241\ : std_logic;
signal \N__1240\ : std_logic;
signal \N__1235\ : std_logic;
signal \N__1232\ : std_logic;
signal \N__1229\ : std_logic;
signal \N__1226\ : std_logic;
signal \N__1225\ : std_logic;
signal \N__1222\ : std_logic;
signal \N__1219\ : std_logic;
signal \N__1216\ : std_logic;
signal \N__1211\ : std_logic;
signal \N__1208\ : std_logic;
signal \N__1205\ : std_logic;
signal \N__1202\ : std_logic;
signal \N__1199\ : std_logic;
signal \N__1196\ : std_logic;
signal \N__1193\ : std_logic;
signal \N__1190\ : std_logic;
signal \N__1187\ : std_logic;
signal \N__1184\ : std_logic;
signal \N__1181\ : std_logic;
signal \N__1180\ : std_logic;
signal \N__1179\ : std_logic;
signal \N__1174\ : std_logic;
signal \N__1171\ : std_logic;
signal \N__1166\ : std_logic;
signal \N__1163\ : std_logic;
signal \N__1160\ : std_logic;
signal \N__1157\ : std_logic;
signal \N__1154\ : std_logic;
signal \N__1151\ : std_logic;
signal \N__1148\ : std_logic;
signal \N__1145\ : std_logic;
signal \N__1142\ : std_logic;
signal \N__1139\ : std_logic;
signal \N__1136\ : std_logic;
signal \N__1133\ : std_logic;
signal \N__1130\ : std_logic;
signal \N__1127\ : std_logic;
signal \N__1124\ : std_logic;
signal \N__1121\ : std_logic;
signal \N__1118\ : std_logic;
signal \N__1115\ : std_logic;
signal \N__1112\ : std_logic;
signal \N__1109\ : std_logic;
signal \N__1106\ : std_logic;
signal \N__1103\ : std_logic;
signal \N__1100\ : std_logic;
signal \N__1097\ : std_logic;
signal \N__1094\ : std_logic;
signal \N__1091\ : std_logic;
signal \N__1090\ : std_logic;
signal \N__1087\ : std_logic;
signal \N__1084\ : std_logic;
signal \N__1079\ : std_logic;
signal \N__1078\ : std_logic;
signal \N__1077\ : std_logic;
signal \N__1076\ : std_logic;
signal \N__1073\ : std_logic;
signal \N__1072\ : std_logic;
signal \N__1071\ : std_logic;
signal \N__1070\ : std_logic;
signal \N__1061\ : std_logic;
signal \N__1058\ : std_logic;
signal \N__1053\ : std_logic;
signal \N__1046\ : std_logic;
signal \N__1045\ : std_logic;
signal \N__1044\ : std_logic;
signal \N__1043\ : std_logic;
signal \N__1040\ : std_logic;
signal \N__1035\ : std_logic;
signal \N__1032\ : std_logic;
signal \N__1025\ : std_logic;
signal \N__1022\ : std_logic;
signal \N__1019\ : std_logic;
signal \N__1016\ : std_logic;
signal \N__1013\ : std_logic;
signal \N__1010\ : std_logic;
signal \N__1007\ : std_logic;
signal \N__1004\ : std_logic;
signal \N__1001\ : std_logic;
signal \N__998\ : std_logic;
signal \N__995\ : std_logic;
signal \N__994\ : std_logic;
signal \N__993\ : std_logic;
signal \N__990\ : std_logic;
signal \N__989\ : std_logic;
signal \N__988\ : std_logic;
signal \N__985\ : std_logic;
signal \N__984\ : std_logic;
signal \N__981\ : std_logic;
signal \N__974\ : std_logic;
signal \N__969\ : std_logic;
signal \N__962\ : std_logic;
signal \N__959\ : std_logic;
signal \N__956\ : std_logic;
signal \N__955\ : std_logic;
signal \N__952\ : std_logic;
signal \N__951\ : std_logic;
signal \N__950\ : std_logic;
signal \N__949\ : std_logic;
signal \N__948\ : std_logic;
signal \N__947\ : std_logic;
signal \N__946\ : std_logic;
signal \N__945\ : std_logic;
signal \N__942\ : std_logic;
signal \N__939\ : std_logic;
signal \N__936\ : std_logic;
signal \N__929\ : std_logic;
signal \N__922\ : std_logic;
signal \N__911\ : std_logic;
signal \N__908\ : std_logic;
signal \N__905\ : std_logic;
signal \N__902\ : std_logic;
signal \N__899\ : std_logic;
signal \N__896\ : std_logic;
signal \N__893\ : std_logic;
signal \N__892\ : std_logic;
signal \N__889\ : std_logic;
signal \N__886\ : std_logic;
signal \N__881\ : std_logic;
signal \N__878\ : std_logic;
signal \N__877\ : std_logic;
signal \N__876\ : std_logic;
signal \N__875\ : std_logic;
signal \N__874\ : std_logic;
signal \N__869\ : std_logic;
signal \N__862\ : std_logic;
signal \N__857\ : std_logic;
signal \N__856\ : std_logic;
signal \N__855\ : std_logic;
signal \N__854\ : std_logic;
signal \N__851\ : std_logic;
signal \N__848\ : std_logic;
signal \N__843\ : std_logic;
signal \N__840\ : std_logic;
signal \N__833\ : std_logic;
signal \N__832\ : std_logic;
signal \N__829\ : std_logic;
signal \N__828\ : std_logic;
signal \N__821\ : std_logic;
signal \N__818\ : std_logic;
signal \N__815\ : std_logic;
signal \N__812\ : std_logic;
signal \N__809\ : std_logic;
signal \N__808\ : std_logic;
signal \N__807\ : std_logic;
signal \N__804\ : std_logic;
signal \N__799\ : std_logic;
signal \N__796\ : std_logic;
signal \N__793\ : std_logic;
signal \N__788\ : std_logic;
signal \N__785\ : std_logic;
signal \N__782\ : std_logic;
signal \N__779\ : std_logic;
signal \N__776\ : std_logic;
signal \N__773\ : std_logic;
signal \N__770\ : std_logic;
signal \N__769\ : std_logic;
signal \N__768\ : std_logic;
signal \N__767\ : std_logic;
signal \N__766\ : std_logic;
signal \N__755\ : std_logic;
signal \N__752\ : std_logic;
signal \N__751\ : std_logic;
signal \N__750\ : std_logic;
signal \N__749\ : std_logic;
signal \N__746\ : std_logic;
signal \N__739\ : std_logic;
signal \N__734\ : std_logic;
signal \N__731\ : std_logic;
signal \N__730\ : std_logic;
signal \N__729\ : std_logic;
signal \N__728\ : std_logic;
signal \N__725\ : std_logic;
signal \N__722\ : std_logic;
signal \N__719\ : std_logic;
signal \N__718\ : std_logic;
signal \N__715\ : std_logic;
signal \N__706\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \RST_N_c_i\ : std_logic;
signal \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.counterZ0Z_0\ : std_logic;
signal \fsm_shiftRegs_inst1.counterZ0Z_1\ : std_logic;
signal \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.counterZ0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.N_123_1\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.counterDYNZ0Z_1\ : std_logic;
signal \fsm_shiftRegs_inst1.counterDYNZ0Z_2\ : std_logic;
signal \fsm_shiftRegs_inst1.counterDYNZ0Z_3\ : std_logic;
signal \RST_N_c\ : std_logic;
signal \fsm_shiftRegs_inst1.current_stateZ0Z_1\ : std_logic;
signal \fsm_shiftRegs_inst1.counterZ0Z_2\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2\ : std_logic;
signal \ENdin_c\ : std_logic;
signal \fsm_shiftRegs_inst1.counterDYNZ0Z_0\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.current_stateZ0Z_2\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_10\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_13\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_14\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_15\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_11\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_12\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_8\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_9\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_6\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_7\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_2\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_4\ : std_logic;
signal \fsm_shiftRegs_inst1.bit_sequenceZ0Z_5\ : std_logic;
signal \fsm_shiftRegs_inst1.un1_current_state4_0\ : std_logic;
signal \fsm_shiftRegs_inst1.current_stateZ0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \fsm_shiftRegs_inst1.current_stateZ0Z_0\ : std_logic;
signal \fsm_shiftRegs_inst1.current_stateZ0Z_4\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0\ : std_logic;
signal \SELSTAT\ : std_logic;
signal signal_out_fsm : std_logic;
signal \SELDYN\ : std_logic;
signal generated_signal_c : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_0\ : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_1\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_0\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_2\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_1\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_3\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_2\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_4\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_3\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_5\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_4\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_6\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_5\ : std_logic;
signal \fsm_shiftRegs_inst1.current_state_i_4\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2_cry_6\ : std_logic;
signal \fsm_shiftRegs_inst1.counter2Z0Z_7\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \CLK_c_g\ : std_logic;
signal \RST_N_c_i_g\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \RST_N_wire\ : std_logic;
signal generated_signal_wire : std_logic;
signal \ENdin_wire\ : std_logic;

begin
    \CLK_wire\ <= CLK;
    \RST_N_wire\ <= RST_N;
    generated_signal <= generated_signal_wire;
    ENdin <= \ENdin_wire\;

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__1626\,
            GLOBALBUFFEROUTPUT => \CLK_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1628\,
            DIN => \N__1627\,
            DOUT => \N__1626\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1628\,
            PADOUT => \N__1627\,
            PADIN => \N__1626\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RST_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1617\,
            DIN => \N__1616\,
            DOUT => \N__1615\,
            PACKAGEPIN => \RST_N_wire\
        );

    \RST_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1617\,
            PADOUT => \N__1616\,
            PADIN => \N__1615\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RST_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \generated_signal_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1608\,
            DIN => \N__1607\,
            DOUT => \N__1606\,
            PACKAGEPIN => generated_signal_wire
        );

    \generated_signal_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1608\,
            PADOUT => \N__1607\,
            PADIN => \N__1606\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1205\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ENdin_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1599\,
            DIN => \N__1598\,
            DOUT => \N__1597\,
            PACKAGEPIN => \ENdin_wire\
        );

    \ENdin_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1599\,
            PADOUT => \N__1598\,
            PADIN => \N__1597\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1016\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__354\ : CascadeMux
    port map (
            O => \N__1580\,
            I => \N__1575\
        );

    \I__353\ : CascadeMux
    port map (
            O => \N__1579\,
            I => \N__1572\
        );

    \I__352\ : CascadeMux
    port map (
            O => \N__1578\,
            I => \N__1569\
        );

    \I__351\ : InMux
    port map (
            O => \N__1575\,
            I => \N__1564\
        );

    \I__350\ : InMux
    port map (
            O => \N__1572\,
            I => \N__1564\
        );

    \I__349\ : InMux
    port map (
            O => \N__1569\,
            I => \N__1561\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__1564\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_1\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__1561\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_1\
        );

    \I__346\ : InMux
    port map (
            O => \N__1556\,
            I => \fsm_shiftRegs_inst1.counter2_cry_0\
        );

    \I__345\ : InMux
    port map (
            O => \N__1553\,
            I => \N__1548\
        );

    \I__344\ : InMux
    port map (
            O => \N__1552\,
            I => \N__1545\
        );

    \I__343\ : InMux
    port map (
            O => \N__1551\,
            I => \N__1542\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__1548\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_2\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__1545\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_2\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__1542\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_2\
        );

    \I__339\ : InMux
    port map (
            O => \N__1535\,
            I => \fsm_shiftRegs_inst1.counter2_cry_1\
        );

    \I__338\ : InMux
    port map (
            O => \N__1532\,
            I => \N__1528\
        );

    \I__337\ : InMux
    port map (
            O => \N__1531\,
            I => \N__1525\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__1528\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_3\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__1525\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_3\
        );

    \I__334\ : InMux
    port map (
            O => \N__1520\,
            I => \fsm_shiftRegs_inst1.counter2_cry_2\
        );

    \I__333\ : CascadeMux
    port map (
            O => \N__1517\,
            I => \N__1512\
        );

    \I__332\ : InMux
    port map (
            O => \N__1516\,
            I => \N__1507\
        );

    \I__331\ : InMux
    port map (
            O => \N__1515\,
            I => \N__1507\
        );

    \I__330\ : InMux
    port map (
            O => \N__1512\,
            I => \N__1504\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__1507\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_4\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__1504\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_4\
        );

    \I__327\ : InMux
    port map (
            O => \N__1499\,
            I => \fsm_shiftRegs_inst1.counter2_cry_3\
        );

    \I__326\ : InMux
    port map (
            O => \N__1496\,
            I => \N__1492\
        );

    \I__325\ : InMux
    port map (
            O => \N__1495\,
            I => \N__1489\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__1492\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_5\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__1489\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_5\
        );

    \I__322\ : InMux
    port map (
            O => \N__1484\,
            I => \fsm_shiftRegs_inst1.counter2_cry_4\
        );

    \I__321\ : CascadeMux
    port map (
            O => \N__1481\,
            I => \N__1478\
        );

    \I__320\ : InMux
    port map (
            O => \N__1478\,
            I => \N__1474\
        );

    \I__319\ : InMux
    port map (
            O => \N__1477\,
            I => \N__1471\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__1474\,
            I => \N__1468\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__1471\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_6\
        );

    \I__316\ : Odrv4
    port map (
            O => \N__1468\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_6\
        );

    \I__315\ : InMux
    port map (
            O => \N__1463\,
            I => \fsm_shiftRegs_inst1.counter2_cry_5\
        );

    \I__314\ : InMux
    port map (
            O => \N__1460\,
            I => \N__1444\
        );

    \I__313\ : InMux
    port map (
            O => \N__1459\,
            I => \N__1444\
        );

    \I__312\ : InMux
    port map (
            O => \N__1458\,
            I => \N__1444\
        );

    \I__311\ : InMux
    port map (
            O => \N__1457\,
            I => \N__1444\
        );

    \I__310\ : InMux
    port map (
            O => \N__1456\,
            I => \N__1435\
        );

    \I__309\ : InMux
    port map (
            O => \N__1455\,
            I => \N__1435\
        );

    \I__308\ : InMux
    port map (
            O => \N__1454\,
            I => \N__1435\
        );

    \I__307\ : InMux
    port map (
            O => \N__1453\,
            I => \N__1435\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__1444\,
            I => \fsm_shiftRegs_inst1.current_state_i_4\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__1435\,
            I => \fsm_shiftRegs_inst1.current_state_i_4\
        );

    \I__304\ : InMux
    port map (
            O => \N__1430\,
            I => \fsm_shiftRegs_inst1.counter2_cry_6\
        );

    \I__303\ : InMux
    port map (
            O => \N__1427\,
            I => \N__1423\
        );

    \I__302\ : InMux
    port map (
            O => \N__1426\,
            I => \N__1420\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__1423\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_7\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__1420\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_7\
        );

    \I__299\ : ClkMux
    port map (
            O => \N__1415\,
            I => \N__1379\
        );

    \I__298\ : ClkMux
    port map (
            O => \N__1414\,
            I => \N__1379\
        );

    \I__297\ : ClkMux
    port map (
            O => \N__1413\,
            I => \N__1379\
        );

    \I__296\ : ClkMux
    port map (
            O => \N__1412\,
            I => \N__1379\
        );

    \I__295\ : ClkMux
    port map (
            O => \N__1411\,
            I => \N__1379\
        );

    \I__294\ : ClkMux
    port map (
            O => \N__1410\,
            I => \N__1379\
        );

    \I__293\ : ClkMux
    port map (
            O => \N__1409\,
            I => \N__1379\
        );

    \I__292\ : ClkMux
    port map (
            O => \N__1408\,
            I => \N__1379\
        );

    \I__291\ : ClkMux
    port map (
            O => \N__1407\,
            I => \N__1379\
        );

    \I__290\ : ClkMux
    port map (
            O => \N__1406\,
            I => \N__1379\
        );

    \I__289\ : ClkMux
    port map (
            O => \N__1405\,
            I => \N__1379\
        );

    \I__288\ : ClkMux
    port map (
            O => \N__1404\,
            I => \N__1379\
        );

    \I__287\ : GlobalMux
    port map (
            O => \N__1379\,
            I => \N__1376\
        );

    \I__286\ : gio2CtrlBuf
    port map (
            O => \N__1376\,
            I => \CLK_c_g\
        );

    \I__285\ : SRMux
    port map (
            O => \N__1373\,
            I => \N__1346\
        );

    \I__284\ : SRMux
    port map (
            O => \N__1372\,
            I => \N__1346\
        );

    \I__283\ : SRMux
    port map (
            O => \N__1371\,
            I => \N__1346\
        );

    \I__282\ : SRMux
    port map (
            O => \N__1370\,
            I => \N__1346\
        );

    \I__281\ : SRMux
    port map (
            O => \N__1369\,
            I => \N__1346\
        );

    \I__280\ : SRMux
    port map (
            O => \N__1368\,
            I => \N__1346\
        );

    \I__279\ : SRMux
    port map (
            O => \N__1367\,
            I => \N__1346\
        );

    \I__278\ : SRMux
    port map (
            O => \N__1366\,
            I => \N__1346\
        );

    \I__277\ : SRMux
    port map (
            O => \N__1365\,
            I => \N__1346\
        );

    \I__276\ : GlobalMux
    port map (
            O => \N__1346\,
            I => \N__1343\
        );

    \I__275\ : gio2CtrlBuf
    port map (
            O => \N__1343\,
            I => \RST_N_c_i_g\
        );

    \I__274\ : InMux
    port map (
            O => \N__1340\,
            I => \N__1336\
        );

    \I__273\ : InMux
    port map (
            O => \N__1339\,
            I => \N__1333\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__1336\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_3\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__1333\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_3\
        );

    \I__270\ : CascadeMux
    port map (
            O => \N__1328\,
            I => \fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_\
        );

    \I__269\ : CascadeMux
    port map (
            O => \N__1325\,
            I => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_\
        );

    \I__268\ : CascadeMux
    port map (
            O => \N__1322\,
            I => \N__1319\
        );

    \I__267\ : InMux
    port map (
            O => \N__1319\,
            I => \N__1316\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__1316\,
            I => \N__1299\
        );

    \I__265\ : InMux
    port map (
            O => \N__1315\,
            I => \N__1286\
        );

    \I__264\ : InMux
    port map (
            O => \N__1314\,
            I => \N__1286\
        );

    \I__263\ : InMux
    port map (
            O => \N__1313\,
            I => \N__1286\
        );

    \I__262\ : InMux
    port map (
            O => \N__1312\,
            I => \N__1286\
        );

    \I__261\ : InMux
    port map (
            O => \N__1311\,
            I => \N__1286\
        );

    \I__260\ : InMux
    port map (
            O => \N__1310\,
            I => \N__1286\
        );

    \I__259\ : InMux
    port map (
            O => \N__1309\,
            I => \N__1269\
        );

    \I__258\ : InMux
    port map (
            O => \N__1308\,
            I => \N__1269\
        );

    \I__257\ : InMux
    port map (
            O => \N__1307\,
            I => \N__1269\
        );

    \I__256\ : InMux
    port map (
            O => \N__1306\,
            I => \N__1269\
        );

    \I__255\ : InMux
    port map (
            O => \N__1305\,
            I => \N__1269\
        );

    \I__254\ : InMux
    port map (
            O => \N__1304\,
            I => \N__1269\
        );

    \I__253\ : InMux
    port map (
            O => \N__1303\,
            I => \N__1269\
        );

    \I__252\ : InMux
    port map (
            O => \N__1302\,
            I => \N__1269\
        );

    \I__251\ : Odrv12
    port map (
            O => \N__1299\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_0\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__1286\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_0\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__1269\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_0\
        );

    \I__248\ : InMux
    port map (
            O => \N__1262\,
            I => \N__1256\
        );

    \I__247\ : InMux
    port map (
            O => \N__1261\,
            I => \N__1253\
        );

    \I__246\ : InMux
    port map (
            O => \N__1260\,
            I => \N__1248\
        );

    \I__245\ : InMux
    port map (
            O => \N__1259\,
            I => \N__1248\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__1256\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_4\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__1253\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_4\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__1248\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_4\
        );

    \I__241\ : InMux
    port map (
            O => \N__1241\,
            I => \N__1235\
        );

    \I__240\ : InMux
    port map (
            O => \N__1240\,
            I => \N__1235\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__1235\,
            I => \fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0\
        );

    \I__238\ : InMux
    port map (
            O => \N__1232\,
            I => \N__1229\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__1229\,
            I => \SELSTAT\
        );

    \I__236\ : InMux
    port map (
            O => \N__1226\,
            I => \N__1222\
        );

    \I__235\ : InMux
    port map (
            O => \N__1225\,
            I => \N__1219\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__1222\,
            I => \N__1216\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__1219\,
            I => signal_out_fsm
        );

    \I__232\ : Odrv12
    port map (
            O => \N__1216\,
            I => signal_out_fsm
        );

    \I__231\ : InMux
    port map (
            O => \N__1211\,
            I => \N__1208\
        );

    \I__230\ : LocalMux
    port map (
            O => \N__1208\,
            I => \SELDYN\
        );

    \I__229\ : IoInMux
    port map (
            O => \N__1205\,
            I => \N__1202\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__1202\,
            I => \N__1199\
        );

    \I__227\ : IoSpan4Mux
    port map (
            O => \N__1199\,
            I => \N__1196\
        );

    \I__226\ : IoSpan4Mux
    port map (
            O => \N__1196\,
            I => \N__1193\
        );

    \I__225\ : Sp12to4
    port map (
            O => \N__1193\,
            I => \N__1190\
        );

    \I__224\ : Span12Mux_s7_h
    port map (
            O => \N__1190\,
            I => \N__1187\
        );

    \I__223\ : Span12Mux_v
    port map (
            O => \N__1187\,
            I => \N__1184\
        );

    \I__222\ : Odrv12
    port map (
            O => \N__1184\,
            I => generated_signal_c
        );

    \I__221\ : InMux
    port map (
            O => \N__1181\,
            I => \N__1174\
        );

    \I__220\ : InMux
    port map (
            O => \N__1180\,
            I => \N__1174\
        );

    \I__219\ : InMux
    port map (
            O => \N__1179\,
            I => \N__1171\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__1174\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_0\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__1171\,
            I => \fsm_shiftRegs_inst1.counter2Z0Z_0\
        );

    \I__216\ : InMux
    port map (
            O => \N__1166\,
            I => \bfn_16_16_0_\
        );

    \I__215\ : InMux
    port map (
            O => \N__1163\,
            I => \N__1160\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__1160\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_14\
        );

    \I__213\ : InMux
    port map (
            O => \N__1157\,
            I => \N__1154\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__1154\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_15\
        );

    \I__211\ : InMux
    port map (
            O => \N__1151\,
            I => \N__1148\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__1148\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_11\
        );

    \I__209\ : InMux
    port map (
            O => \N__1145\,
            I => \N__1142\
        );

    \I__208\ : LocalMux
    port map (
            O => \N__1142\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_12\
        );

    \I__207\ : InMux
    port map (
            O => \N__1139\,
            I => \N__1136\
        );

    \I__206\ : LocalMux
    port map (
            O => \N__1136\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_8\
        );

    \I__205\ : InMux
    port map (
            O => \N__1133\,
            I => \N__1130\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__1130\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_9\
        );

    \I__203\ : InMux
    port map (
            O => \N__1127\,
            I => \N__1124\
        );

    \I__202\ : LocalMux
    port map (
            O => \N__1124\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_6\
        );

    \I__201\ : InMux
    port map (
            O => \N__1121\,
            I => \N__1118\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__1118\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_7\
        );

    \I__199\ : InMux
    port map (
            O => \N__1115\,
            I => \N__1112\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__1112\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_2\
        );

    \I__197\ : InMux
    port map (
            O => \N__1109\,
            I => \N__1106\
        );

    \I__196\ : LocalMux
    port map (
            O => \N__1106\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_3\
        );

    \I__195\ : InMux
    port map (
            O => \N__1103\,
            I => \N__1100\
        );

    \I__194\ : LocalMux
    port map (
            O => \N__1100\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_4\
        );

    \I__193\ : InMux
    port map (
            O => \N__1097\,
            I => \N__1094\
        );

    \I__192\ : LocalMux
    port map (
            O => \N__1094\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_5\
        );

    \I__191\ : CEMux
    port map (
            O => \N__1091\,
            I => \N__1087\
        );

    \I__190\ : CEMux
    port map (
            O => \N__1090\,
            I => \N__1084\
        );

    \I__189\ : LocalMux
    port map (
            O => \N__1087\,
            I => \fsm_shiftRegs_inst1.un1_current_state4_0\
        );

    \I__188\ : LocalMux
    port map (
            O => \N__1084\,
            I => \fsm_shiftRegs_inst1.un1_current_state4_0\
        );

    \I__187\ : CascadeMux
    port map (
            O => \N__1079\,
            I => \N__1073\
        );

    \I__186\ : InMux
    port map (
            O => \N__1078\,
            I => \N__1061\
        );

    \I__185\ : InMux
    port map (
            O => \N__1077\,
            I => \N__1061\
        );

    \I__184\ : InMux
    port map (
            O => \N__1076\,
            I => \N__1061\
        );

    \I__183\ : InMux
    port map (
            O => \N__1073\,
            I => \N__1061\
        );

    \I__182\ : InMux
    port map (
            O => \N__1072\,
            I => \N__1058\
        );

    \I__181\ : InMux
    port map (
            O => \N__1071\,
            I => \N__1053\
        );

    \I__180\ : InMux
    port map (
            O => \N__1070\,
            I => \N__1053\
        );

    \I__179\ : LocalMux
    port map (
            O => \N__1061\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_1\
        );

    \I__178\ : LocalMux
    port map (
            O => \N__1058\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_1\
        );

    \I__177\ : LocalMux
    port map (
            O => \N__1053\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_1\
        );

    \I__176\ : InMux
    port map (
            O => \N__1046\,
            I => \N__1040\
        );

    \I__175\ : InMux
    port map (
            O => \N__1045\,
            I => \N__1035\
        );

    \I__174\ : InMux
    port map (
            O => \N__1044\,
            I => \N__1035\
        );

    \I__173\ : InMux
    port map (
            O => \N__1043\,
            I => \N__1032\
        );

    \I__172\ : LocalMux
    port map (
            O => \N__1040\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_2\
        );

    \I__171\ : LocalMux
    port map (
            O => \N__1035\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_2\
        );

    \I__170\ : LocalMux
    port map (
            O => \N__1032\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_2\
        );

    \I__169\ : InMux
    port map (
            O => \N__1025\,
            I => \N__1022\
        );

    \I__168\ : LocalMux
    port map (
            O => \N__1022\,
            I => \N__1019\
        );

    \I__167\ : Odrv4
    port map (
            O => \N__1019\,
            I => \fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2\
        );

    \I__166\ : IoInMux
    port map (
            O => \N__1016\,
            I => \N__1013\
        );

    \I__165\ : LocalMux
    port map (
            O => \N__1013\,
            I => \N__1010\
        );

    \I__164\ : IoSpan4Mux
    port map (
            O => \N__1010\,
            I => \N__1007\
        );

    \I__163\ : Span4Mux_s3_h
    port map (
            O => \N__1007\,
            I => \N__1004\
        );

    \I__162\ : Sp12to4
    port map (
            O => \N__1004\,
            I => \N__1001\
        );

    \I__161\ : Span12Mux_h
    port map (
            O => \N__1001\,
            I => \N__998\
        );

    \I__160\ : Odrv12
    port map (
            O => \N__998\,
            I => \ENdin_c\
        );

    \I__159\ : CascadeMux
    port map (
            O => \N__995\,
            I => \N__990\
        );

    \I__158\ : CascadeMux
    port map (
            O => \N__994\,
            I => \N__985\
        );

    \I__157\ : InMux
    port map (
            O => \N__993\,
            I => \N__981\
        );

    \I__156\ : InMux
    port map (
            O => \N__990\,
            I => \N__974\
        );

    \I__155\ : InMux
    port map (
            O => \N__989\,
            I => \N__974\
        );

    \I__154\ : InMux
    port map (
            O => \N__988\,
            I => \N__974\
        );

    \I__153\ : InMux
    port map (
            O => \N__985\,
            I => \N__969\
        );

    \I__152\ : InMux
    port map (
            O => \N__984\,
            I => \N__969\
        );

    \I__151\ : LocalMux
    port map (
            O => \N__981\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_0\
        );

    \I__150\ : LocalMux
    port map (
            O => \N__974\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_0\
        );

    \I__149\ : LocalMux
    port map (
            O => \N__969\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_0\
        );

    \I__148\ : InMux
    port map (
            O => \N__962\,
            I => \N__959\
        );

    \I__147\ : LocalMux
    port map (
            O => \N__959\,
            I => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3\
        );

    \I__146\ : CascadeMux
    port map (
            O => \N__956\,
            I => \N__952\
        );

    \I__145\ : InMux
    port map (
            O => \N__955\,
            I => \N__942\
        );

    \I__144\ : InMux
    port map (
            O => \N__952\,
            I => \N__939\
        );

    \I__143\ : InMux
    port map (
            O => \N__951\,
            I => \N__936\
        );

    \I__142\ : InMux
    port map (
            O => \N__950\,
            I => \N__929\
        );

    \I__141\ : InMux
    port map (
            O => \N__949\,
            I => \N__929\
        );

    \I__140\ : InMux
    port map (
            O => \N__948\,
            I => \N__929\
        );

    \I__139\ : InMux
    port map (
            O => \N__947\,
            I => \N__922\
        );

    \I__138\ : InMux
    port map (
            O => \N__946\,
            I => \N__922\
        );

    \I__137\ : InMux
    port map (
            O => \N__945\,
            I => \N__922\
        );

    \I__136\ : LocalMux
    port map (
            O => \N__942\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_2\
        );

    \I__135\ : LocalMux
    port map (
            O => \N__939\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_2\
        );

    \I__134\ : LocalMux
    port map (
            O => \N__936\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_2\
        );

    \I__133\ : LocalMux
    port map (
            O => \N__929\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_2\
        );

    \I__132\ : LocalMux
    port map (
            O => \N__922\,
            I => \fsm_shiftRegs_inst1.current_stateZ0Z_2\
        );

    \I__131\ : InMux
    port map (
            O => \N__911\,
            I => \N__908\
        );

    \I__130\ : LocalMux
    port map (
            O => \N__908\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_10\
        );

    \I__129\ : InMux
    port map (
            O => \N__905\,
            I => \N__902\
        );

    \I__128\ : LocalMux
    port map (
            O => \N__902\,
            I => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_13\
        );

    \I__127\ : CascadeMux
    port map (
            O => \N__899\,
            I => \fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_\
        );

    \I__126\ : InMux
    port map (
            O => \N__896\,
            I => \N__893\
        );

    \I__125\ : LocalMux
    port map (
            O => \N__893\,
            I => \N__889\
        );

    \I__124\ : InMux
    port map (
            O => \N__892\,
            I => \N__886\
        );

    \I__123\ : Odrv4
    port map (
            O => \N__889\,
            I => \fsm_shiftRegs_inst1.N_123_1\
        );

    \I__122\ : LocalMux
    port map (
            O => \N__886\,
            I => \fsm_shiftRegs_inst1.N_123_1\
        );

    \I__121\ : CascadeMux
    port map (
            O => \N__881\,
            I => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_\
        );

    \I__120\ : InMux
    port map (
            O => \N__878\,
            I => \N__869\
        );

    \I__119\ : InMux
    port map (
            O => \N__877\,
            I => \N__869\
        );

    \I__118\ : InMux
    port map (
            O => \N__876\,
            I => \N__862\
        );

    \I__117\ : InMux
    port map (
            O => \N__875\,
            I => \N__862\
        );

    \I__116\ : InMux
    port map (
            O => \N__874\,
            I => \N__862\
        );

    \I__115\ : LocalMux
    port map (
            O => \N__869\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_1\
        );

    \I__114\ : LocalMux
    port map (
            O => \N__862\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_1\
        );

    \I__113\ : CascadeMux
    port map (
            O => \N__857\,
            I => \N__851\
        );

    \I__112\ : InMux
    port map (
            O => \N__856\,
            I => \N__848\
        );

    \I__111\ : InMux
    port map (
            O => \N__855\,
            I => \N__843\
        );

    \I__110\ : InMux
    port map (
            O => \N__854\,
            I => \N__843\
        );

    \I__109\ : InMux
    port map (
            O => \N__851\,
            I => \N__840\
        );

    \I__108\ : LocalMux
    port map (
            O => \N__848\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_2\
        );

    \I__107\ : LocalMux
    port map (
            O => \N__843\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_2\
        );

    \I__106\ : LocalMux
    port map (
            O => \N__840\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_2\
        );

    \I__105\ : CascadeMux
    port map (
            O => \N__833\,
            I => \N__829\
        );

    \I__104\ : InMux
    port map (
            O => \N__832\,
            I => \N__821\
        );

    \I__103\ : InMux
    port map (
            O => \N__829\,
            I => \N__821\
        );

    \I__102\ : InMux
    port map (
            O => \N__828\,
            I => \N__821\
        );

    \I__101\ : LocalMux
    port map (
            O => \N__821\,
            I => \fsm_shiftRegs_inst1.counterDYNZ0Z_3\
        );

    \I__100\ : InMux
    port map (
            O => \N__818\,
            I => \N__815\
        );

    \I__99\ : LocalMux
    port map (
            O => \N__815\,
            I => \N__812\
        );

    \I__98\ : Span4Mux_v
    port map (
            O => \N__812\,
            I => \N__809\
        );

    \I__97\ : Span4Mux_v
    port map (
            O => \N__809\,
            I => \N__804\
        );

    \I__96\ : InMux
    port map (
            O => \N__808\,
            I => \N__799\
        );

    \I__95\ : InMux
    port map (
            O => \N__807\,
            I => \N__799\
        );

    \I__94\ : Sp12to4
    port map (
            O => \N__804\,
            I => \N__796\
        );

    \I__93\ : LocalMux
    port map (
            O => \N__799\,
            I => \N__793\
        );

    \I__92\ : Span12Mux_h
    port map (
            O => \N__796\,
            I => \N__788\
        );

    \I__91\ : Span12Mux_v
    port map (
            O => \N__793\,
            I => \N__788\
        );

    \I__90\ : Span12Mux_h
    port map (
            O => \N__788\,
            I => \N__785\
        );

    \I__89\ : Odrv12
    port map (
            O => \N__785\,
            I => \RST_N_c\
        );

    \I__88\ : IoInMux
    port map (
            O => \N__782\,
            I => \N__779\
        );

    \I__87\ : LocalMux
    port map (
            O => \N__779\,
            I => \N__776\
        );

    \I__86\ : Odrv12
    port map (
            O => \N__776\,
            I => \RST_N_c_i\
        );

    \I__85\ : CascadeMux
    port map (
            O => \N__773\,
            I => \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_\
        );

    \I__84\ : InMux
    port map (
            O => \N__770\,
            I => \N__755\
        );

    \I__83\ : InMux
    port map (
            O => \N__769\,
            I => \N__755\
        );

    \I__82\ : InMux
    port map (
            O => \N__768\,
            I => \N__755\
        );

    \I__81\ : InMux
    port map (
            O => \N__767\,
            I => \N__755\
        );

    \I__80\ : InMux
    port map (
            O => \N__766\,
            I => \N__755\
        );

    \I__79\ : LocalMux
    port map (
            O => \N__755\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_0\
        );

    \I__78\ : InMux
    port map (
            O => \N__752\,
            I => \N__746\
        );

    \I__77\ : InMux
    port map (
            O => \N__751\,
            I => \N__739\
        );

    \I__76\ : InMux
    port map (
            O => \N__750\,
            I => \N__739\
        );

    \I__75\ : InMux
    port map (
            O => \N__749\,
            I => \N__739\
        );

    \I__74\ : LocalMux
    port map (
            O => \N__746\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_1\
        );

    \I__73\ : LocalMux
    port map (
            O => \N__739\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_1\
        );

    \I__72\ : CascadeMux
    port map (
            O => \N__734\,
            I => \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3_cascade_\
        );

    \I__71\ : CascadeMux
    port map (
            O => \N__731\,
            I => \N__725\
        );

    \I__70\ : CascadeMux
    port map (
            O => \N__730\,
            I => \N__722\
        );

    \I__69\ : CascadeMux
    port map (
            O => \N__729\,
            I => \N__719\
        );

    \I__68\ : InMux
    port map (
            O => \N__728\,
            I => \N__715\
        );

    \I__67\ : InMux
    port map (
            O => \N__725\,
            I => \N__706\
        );

    \I__66\ : InMux
    port map (
            O => \N__722\,
            I => \N__706\
        );

    \I__65\ : InMux
    port map (
            O => \N__719\,
            I => \N__706\
        );

    \I__64\ : InMux
    port map (
            O => \N__718\,
            I => \N__706\
        );

    \I__63\ : LocalMux
    port map (
            O => \N__715\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_3\
        );

    \I__62\ : LocalMux
    port map (
            O => \N__706\,
            I => \fsm_shiftRegs_inst1.counterZ0Z_3\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_16_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \RST_N_ibuf_RNIBJGC_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__782\,
            GLOBALBUFFEROUTPUT => \RST_N_c_i_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \RST_N_ibuf_RNIBJGC_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__818\,
            lcout => \RST_N_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counter_RNO_0_2_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100001000"
        )
    port map (
            in0 => \N__767\,
            in1 => \N__750\,
            in2 => \N__729\,
            in3 => \N__1044\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counter_2_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__1076\,
            in1 => \_gnd_net_\,
            in2 => \N__773\,
            in3 => \_gnd_net_\,
            lcout => \fsm_shiftRegs_inst1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1405\,
            ce => 'H',
            sr => \N__1366\
        );

    \fsm_shiftRegs_inst1.counter_0_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010100000000"
        )
    port map (
            in0 => \N__769\,
            in1 => \_gnd_net_\,
            in2 => \N__731\,
            in3 => \N__1078\,
            lcout => \fsm_shiftRegs_inst1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1405\,
            ce => 'H',
            sr => \N__1366\
        );

    \fsm_shiftRegs_inst1.counter_RNIC589_1_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__749\,
            in1 => \N__766\,
            in2 => \_gnd_net_\,
            in3 => \N__718\,
            lcout => \fsm_shiftRegs_inst1.N_123_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counter_1_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001000011000000"
        )
    port map (
            in0 => \N__728\,
            in1 => \N__752\,
            in2 => \N__1079\,
            in3 => \N__770\,
            lcout => \fsm_shiftRegs_inst1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1405\,
            ce => 'H',
            sr => \N__1366\
        );

    \fsm_shiftRegs_inst1.counter_RNO_0_3_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__768\,
            in1 => \N__751\,
            in2 => \N__730\,
            in3 => \N__1045\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.counter_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counter_3_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__1077\,
            in1 => \_gnd_net_\,
            in2 => \N__734\,
            in3 => \_gnd_net_\,
            lcout => \fsm_shiftRegs_inst1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1405\,
            ce => 'H',
            sr => \N__1366\
        );

    \fsm_shiftRegs_inst1.current_state_1_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011111010"
        )
    port map (
            in0 => \N__1072\,
            in1 => \N__1046\,
            in2 => \N__1322\,
            in3 => \N__892\,
            lcout => \fsm_shiftRegs_inst1.current_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1404\,
            ce => 'H',
            sr => \N__1365\
        );

    \fsm_shiftRegs_inst1.counterDYN_1_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__948\,
            in1 => \N__989\,
            in2 => \_gnd_net_\,
            in3 => \N__878\,
            lcout => \fsm_shiftRegs_inst1.counterDYNZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1411\,
            ce => 'H',
            sr => \N__1369\
        );

    \fsm_shiftRegs_inst1.counterDYN_2_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100110010000000"
        )
    port map (
            in0 => \N__877\,
            in1 => \N__950\,
            in2 => \N__995\,
            in3 => \N__856\,
            lcout => \fsm_shiftRegs_inst1.counterDYNZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1411\,
            ce => 'H',
            sr => \N__1369\
        );

    \fsm_shiftRegs_inst1.counterDYN_0_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__949\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__988\,
            lcout => \fsm_shiftRegs_inst1.counterDYNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1411\,
            ce => 'H',
            sr => \N__1369\
        );

    \fsm_shiftRegs_inst1.counterDYN_RNO_0_3_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__854\,
            in1 => \N__875\,
            in2 => \N__833\,
            in3 => \N__984\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.counterDYN_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counterDYN_3_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__899\,
            in3 => \N__947\,
            lcout => \fsm_shiftRegs_inst1.counterDYNZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1408\,
            ce => 'H',
            sr => \N__1368\
        );

    \fsm_shiftRegs_inst1.current_state_RNO_0_2_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__876\,
            in1 => \N__855\,
            in2 => \N__994\,
            in3 => \N__832\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_2_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__946\,
            in1 => \N__896\,
            in2 => \N__881\,
            in3 => \N__1025\,
            lcout => \fsm_shiftRegs_inst1.current_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1408\,
            ce => 'H',
            sr => \N__1368\
        );

    \fsm_shiftRegs_inst1.current_state_RNO_0_3_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__874\,
            in1 => \N__945\,
            in2 => \N__857\,
            in3 => \N__828\,
            lcout => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.signal_out_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__1225\,
            in1 => \N__1157\,
            in2 => \N__956\,
            in3 => \N__808\,
            lcout => signal_out_fsm,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_RNI7RPG_1_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1070\,
            in2 => \_gnd_net_\,
            in3 => \N__807\,
            lcout => \fsm_shiftRegs_inst1.un1_current_state4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_RNO_1_2_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__1071\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1043\,
            lcout => \fsm_shiftRegs_inst1.current_state_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.en_fin_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__955\,
            lcout => \ENdin_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1414\,
            ce => 'H',
            sr => \N__1372\
        );

    \fsm_shiftRegs_inst1.current_state_3_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__993\,
            in2 => \_gnd_net_\,
            in3 => \N__962\,
            lcout => \fsm_shiftRegs_inst1.current_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1412\,
            ce => 'H',
            sr => \N__1370\
        );

    \fsm_shiftRegs_inst1.sel_dyn_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__951\,
            in2 => \_gnd_net_\,
            in3 => \N__1262\,
            lcout => \SELDYN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1412\,
            ce => 'H',
            sr => \N__1370\
        );

    \fsm_shiftRegs_inst1.bit_sequence_10_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1302\,
            in2 => \_gnd_net_\,
            in3 => \N__1133\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1409\,
            ce => \N__1090\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_11_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__1303\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__911\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1409\,
            ce => \N__1090\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_13_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1305\,
            in2 => \_gnd_net_\,
            in3 => \N__1145\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1409\,
            ce => \N__1090\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_14_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__1306\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__905\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1409\,
            ce => \N__1090\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_8_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1308\,
            in2 => \_gnd_net_\,
            in3 => \N__1121\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1409\,
            ce => \N__1090\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_15_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__1307\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1163\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1409\,
            ce => \N__1090\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_12_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1304\,
            in2 => \_gnd_net_\,
            in3 => \N__1151\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1409\,
            ce => \N__1090\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_9_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__1309\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1139\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1409\,
            ce => \N__1090\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_6_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1313\,
            in2 => \_gnd_net_\,
            in3 => \N__1097\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1407\,
            ce => \N__1091\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_2_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__1315\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1407\,
            ce => \N__1091\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_7_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__1314\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1127\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1407\,
            ce => \N__1091\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_3_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1310\,
            in2 => \_gnd_net_\,
            in3 => \N__1115\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1407\,
            ce => \N__1091\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_4_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__1311\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1109\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1407\,
            ce => \N__1091\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.bit_sequence_5_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1312\,
            in2 => \_gnd_net_\,
            in3 => \N__1103\,
            lcout => \fsm_shiftRegs_inst1.bit_sequenceZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1407\,
            ce => \N__1091\,
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.sel_stat_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1340\,
            lcout => \SELSTAT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1415\,
            ce => 'H',
            sr => \N__1373\
        );

    \fsm_shiftRegs_inst1.current_state_RNO_0_4_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__1553\,
            in1 => \N__1180\,
            in2 => \N__1580\,
            in3 => \N__1516\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.current_state_ns_a3_7_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_4_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111011101110"
        )
    port map (
            in0 => \N__1260\,
            in1 => \N__1339\,
            in2 => \N__1328\,
            in3 => \N__1241\,
            lcout => \fsm_shiftRegs_inst1.current_stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1413\,
            ce => 'H',
            sr => \N__1371\
        );

    \fsm_shiftRegs_inst1.current_state_RNO_0_0_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1552\,
            in2 => \N__1579\,
            in3 => \N__1515\,
            lcout => OPEN,
            ltout => \fsm_shiftRegs_inst1.current_state_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.current_state_0_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__1181\,
            in1 => \N__1261\,
            in2 => \N__1325\,
            in3 => \N__1240\,
            lcout => \fsm_shiftRegs_inst1.current_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1413\,
            ce => 'H',
            sr => \N__1371\
        );

    \fsm_shiftRegs_inst1.current_state_RNIVA94_4_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1259\,
            lcout => \fsm_shiftRegs_inst1.current_state_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_shiftRegs_inst1.counter2_RNITAO81_7_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1495\,
            in1 => \N__1531\,
            in2 => \N__1481\,
            in3 => \N__1426\,
            lcout => \fsm_shiftRegs_inst1.current_state_ns_a3_7_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generator_inst1.signal_aux_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__1232\,
            in1 => \N__1226\,
            in2 => \_gnd_net_\,
            in3 => \N__1211\,
            lcout => generated_signal_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1413\,
            ce => 'H',
            sr => \N__1371\
        );

    \fsm_shiftRegs_inst1.counter2_0_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1457\,
            in1 => \N__1179\,
            in2 => \_gnd_net_\,
            in3 => \N__1166\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_16_16_0_\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_0\,
            clk => \N__1410\,
            ce => 'H',
            sr => \N__1367\
        );

    \fsm_shiftRegs_inst1.counter2_1_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__1453\,
            in1 => \_gnd_net_\,
            in2 => \N__1578\,
            in3 => \N__1556\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_1\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_0\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_1\,
            clk => \N__1410\,
            ce => 'H',
            sr => \N__1367\
        );

    \fsm_shiftRegs_inst1.counter2_2_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1458\,
            in1 => \N__1551\,
            in2 => \_gnd_net_\,
            in3 => \N__1535\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_2\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_1\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_2\,
            clk => \N__1410\,
            ce => 'H',
            sr => \N__1367\
        );

    \fsm_shiftRegs_inst1.counter2_3_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1454\,
            in1 => \N__1532\,
            in2 => \_gnd_net_\,
            in3 => \N__1520\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_3\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_2\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_3\,
            clk => \N__1410\,
            ce => 'H',
            sr => \N__1367\
        );

    \fsm_shiftRegs_inst1.counter2_4_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__1459\,
            in1 => \_gnd_net_\,
            in2 => \N__1517\,
            in3 => \N__1499\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_4\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_3\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_4\,
            clk => \N__1410\,
            ce => 'H',
            sr => \N__1367\
        );

    \fsm_shiftRegs_inst1.counter2_5_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1455\,
            in1 => \N__1496\,
            in2 => \_gnd_net_\,
            in3 => \N__1484\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_5\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_4\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_5\,
            clk => \N__1410\,
            ce => 'H',
            sr => \N__1367\
        );

    \fsm_shiftRegs_inst1.counter2_6_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1460\,
            in1 => \N__1477\,
            in2 => \_gnd_net_\,
            in3 => \N__1463\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_6\,
            ltout => OPEN,
            carryin => \fsm_shiftRegs_inst1.counter2_cry_5\,
            carryout => \fsm_shiftRegs_inst1.counter2_cry_6\,
            clk => \N__1410\,
            ce => 'H',
            sr => \N__1367\
        );

    \fsm_shiftRegs_inst1.counter2_7_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1456\,
            in1 => \N__1427\,
            in2 => \_gnd_net_\,
            in3 => \N__1430\,
            lcout => \fsm_shiftRegs_inst1.counter2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1410\,
            ce => 'H',
            sr => \N__1367\
        );
end \INTERFACE\;
