-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 19 2025 17:18:55

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    SDO_signal_out : out std_logic;
    RST_N : in std_logic;
    CLK : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__5865\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3507\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3333\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3303\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3219\ : std_logic;
signal \N__3216\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3144\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3021\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2997\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \RST_N_c\ : std_logic;
signal \RST_N_c_i\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_72\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_71\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_64\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_65\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_73\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_74\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_75\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_35\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_79\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_78\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_76\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_77\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_34\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_33\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_80\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_81\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_2\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_70\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_68\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_69\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_66\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_67\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_14\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_15\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_13\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_63\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_40\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_41\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_12\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_39\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_36\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_37\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_38\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_1\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_11\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_62\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_60\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_61\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_82\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_32\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_10\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_9\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_31\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_3\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_4\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_59\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_30\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_8\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_29\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_25\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_26\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_5\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_6\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_7\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_27\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_28\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_58\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_16\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_42\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_19\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_17\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_18\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_20\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_21\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_22\ : std_logic;
signal \bfn_3_18_0_\ : std_logic;
signal \fsm_ctrl_inst1.counter_stat_cry_0\ : std_logic;
signal \fsm_ctrl_inst1.counter_stat_cry_1\ : std_logic;
signal \fsm_ctrl_inst1.counter_stat_cry_2\ : std_logic;
signal \fsm_ctrl_inst1.counter_stat_cry_3\ : std_logic;
signal \fsm_ctrl_inst1.counter_stat_cry_4\ : std_logic;
signal \fsm_ctrl_inst1.counter_stat_cry_5\ : std_logic;
signal \fsm_ctrl_inst1.current_state_ns_0_i_0_1_0_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.counter_statZ0Z_1\ : std_logic;
signal \fsm_ctrl_inst1.counter_statZ0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.counter_statZ0Z_2\ : std_logic;
signal \fsm_ctrl_inst1.current_state_ns_i_i_a2_0_4_1_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.current_state_ns_i_i_a2_0_5_1_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.current_state_i_0\ : std_logic;
signal \fsm_ctrl_inst1.counter_idleZ0Z_0\ : std_logic;
signal \bfn_3_20_0_\ : std_logic;
signal \fsm_ctrl_inst1.counter_idleZ0Z_1\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_cry_0\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_cry_1\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_cry_2\ : std_logic;
signal \fsm_ctrl_inst1.counter_idle_cry_3\ : std_logic;
signal \fsm_ctrl_inst1.counter_idlee_0_i\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_56\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_57\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_54\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_55\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_23\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_24\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_48\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_49\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_45\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_43\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_44\ : std_logic;
signal \fsm_ctrl_inst1.counter_statZ0Z_4\ : std_logic;
signal \fsm_ctrl_inst1.counter_statZ0Z_3\ : std_logic;
signal \fsm_ctrl_inst1.counter_statZ0Z_5\ : std_logic;
signal \fsm_ctrl_inst1.counter_statZ0Z_6\ : std_logic;
signal \fsm_ctrl_inst1.counter_stat_RNIML9Z0Z_6_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.counter_stat12_i_0\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_1\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_2\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_3\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_4\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_5\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_6\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_7\ : std_logic;
signal \fsm_ctrl_inst1.counter_state_0_i\ : std_logic;
signal \fsm_ctrl_inst1.counter_idleZ0Z_3\ : std_logic;
signal \fsm_ctrl_inst1.counter_idleZ0Z_2\ : std_logic;
signal \fsm_ctrl_inst1.counter_idleZ0Z_4\ : std_logic;
signal \fsm_ctrl_inst1.N_127_1\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_10\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_11\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_12\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_13\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_14\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_8\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_9\ : std_logic;
signal \fsm_ctrl_inst1.current_state_i_1\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_46\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_47\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_53\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_52\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_50\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_51\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_83\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_84\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_85\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_86\ : std_logic;
signal \fsm_ctrl_inst1.current_state_i_g_0\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_dinZ0Z_15\ : std_logic;
signal \fsm_ctrl_inst1.bit_sequence_statZ0Z_87\ : std_logic;
signal \fsm_ctrl_inst1.current_stateZ0Z_1\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_1\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_0\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_2\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_3\ : std_logic;
signal \MOSI\ : std_logic;
signal \SDO_signal_out_c\ : std_logic;
signal \fsm_ctrl_inst1.counter_din_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \fsm_ctrl_inst1.counter_dinZ0Z_3\ : std_logic;
signal \fsm_ctrl_inst1.counter_din_RNI6L3H1Z0Z_3\ : std_logic;
signal \fsm_ctrl_inst1.counter_dinZ0Z_2\ : std_logic;
signal \fsm_ctrl_inst1.counter_dinZ0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.counter_dinZ0Z_1\ : std_logic;
signal \fsm_ctrl_inst1.current_stateZ0Z_0\ : std_logic;
signal \fsm_ctrl_inst1.SEL_REG_i\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_4\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_5\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_6\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_0\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_1\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_2\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_3\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_12\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_15\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_13\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_14\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_7\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_8\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_9\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_10\ : std_logic;
signal \config_register_latched_dec_inst1.DYNSRZ0Z_11\ : std_logic;
signal \SEL_REG\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_4\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_5\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_6\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_7\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_10\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_8\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_9\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_11\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_12\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_13\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_14\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_15\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_86\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_87\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_85\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_84\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_83\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_16\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_82\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_81\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_17\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_80\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_33\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_32\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_27\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_30\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_31\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_28\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_29\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_25\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_26\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_34\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_23\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_24\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_79\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_18\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_78\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_21\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_22\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_19\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_20\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_75\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_76\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_77\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_73\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_74\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_71\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_72\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_35\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_36\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_37\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_38\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_70\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_66\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_67\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_68\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_69\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_39\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_40\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_41\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_42\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_43\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_59\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_60\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_57\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_58\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_61\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_62\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_63\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_64\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_65\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_46\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_44\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_45\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_47\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_48\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_49\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_50\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_51\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_52\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_53\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_56\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_54\ : std_logic;
signal \config_register_latched_dec_inst1.STATSRZ0Z_55\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \CLK_c_g\ : std_logic;
signal \SEL_REG_i_g\ : std_logic;
signal \RST_N_c_i_g\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \RST_N_wire\ : std_logic;
signal \SDO_signal_out_wire\ : std_logic;

begin
    \CLK_wire\ <= CLK;
    \RST_N_wire\ <= RST_N;
    SDO_signal_out <= \SDO_signal_out_wire\;

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__5863\,
            GLOBALBUFFEROUTPUT => \CLK_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5865\,
            DIN => \N__5864\,
            DOUT => \N__5863\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5865\,
            PADOUT => \N__5864\,
            PADIN => \N__5863\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RST_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5854\,
            DIN => \N__5853\,
            DOUT => \N__5852\,
            PACKAGEPIN => \RST_N_wire\
        );

    \RST_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5854\,
            PADOUT => \N__5853\,
            PADIN => \N__5852\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RST_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SDO_signal_out_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5845\,
            DIN => \N__5844\,
            DOUT => \N__5843\,
            PACKAGEPIN => \SDO_signal_out_wire\
        );

    \SDO_signal_out_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__5845\,
            PADOUT => \N__5844\,
            PADIN => \N__5843\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4542\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1198\ : InMux
    port map (
            O => \N__5826\,
            I => \N__5823\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5823\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_47\
        );

    \I__1196\ : InMux
    port map (
            O => \N__5820\,
            I => \N__5817\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__5817\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_48\
        );

    \I__1194\ : InMux
    port map (
            O => \N__5814\,
            I => \N__5811\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__5811\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_49\
        );

    \I__1192\ : InMux
    port map (
            O => \N__5808\,
            I => \N__5805\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__5805\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_50\
        );

    \I__1190\ : InMux
    port map (
            O => \N__5802\,
            I => \N__5799\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5799\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_51\
        );

    \I__1188\ : InMux
    port map (
            O => \N__5796\,
            I => \N__5793\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5793\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_52\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5790\,
            I => \N__5787\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__5787\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_53\
        );

    \I__1184\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5781\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__5781\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_56\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5778\,
            I => \N__5775\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5775\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_54\
        );

    \I__1180\ : InMux
    port map (
            O => \N__5772\,
            I => \N__5769\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__5769\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_55\
        );

    \I__1178\ : ClkMux
    port map (
            O => \N__5766\,
            I => \N__5595\
        );

    \I__1177\ : ClkMux
    port map (
            O => \N__5765\,
            I => \N__5595\
        );

    \I__1176\ : ClkMux
    port map (
            O => \N__5764\,
            I => \N__5595\
        );

    \I__1175\ : ClkMux
    port map (
            O => \N__5763\,
            I => \N__5595\
        );

    \I__1174\ : ClkMux
    port map (
            O => \N__5762\,
            I => \N__5595\
        );

    \I__1173\ : ClkMux
    port map (
            O => \N__5761\,
            I => \N__5595\
        );

    \I__1172\ : ClkMux
    port map (
            O => \N__5760\,
            I => \N__5595\
        );

    \I__1171\ : ClkMux
    port map (
            O => \N__5759\,
            I => \N__5595\
        );

    \I__1170\ : ClkMux
    port map (
            O => \N__5758\,
            I => \N__5595\
        );

    \I__1169\ : ClkMux
    port map (
            O => \N__5757\,
            I => \N__5595\
        );

    \I__1168\ : ClkMux
    port map (
            O => \N__5756\,
            I => \N__5595\
        );

    \I__1167\ : ClkMux
    port map (
            O => \N__5755\,
            I => \N__5595\
        );

    \I__1166\ : ClkMux
    port map (
            O => \N__5754\,
            I => \N__5595\
        );

    \I__1165\ : ClkMux
    port map (
            O => \N__5753\,
            I => \N__5595\
        );

    \I__1164\ : ClkMux
    port map (
            O => \N__5752\,
            I => \N__5595\
        );

    \I__1163\ : ClkMux
    port map (
            O => \N__5751\,
            I => \N__5595\
        );

    \I__1162\ : ClkMux
    port map (
            O => \N__5750\,
            I => \N__5595\
        );

    \I__1161\ : ClkMux
    port map (
            O => \N__5749\,
            I => \N__5595\
        );

    \I__1160\ : ClkMux
    port map (
            O => \N__5748\,
            I => \N__5595\
        );

    \I__1159\ : ClkMux
    port map (
            O => \N__5747\,
            I => \N__5595\
        );

    \I__1158\ : ClkMux
    port map (
            O => \N__5746\,
            I => \N__5595\
        );

    \I__1157\ : ClkMux
    port map (
            O => \N__5745\,
            I => \N__5595\
        );

    \I__1156\ : ClkMux
    port map (
            O => \N__5744\,
            I => \N__5595\
        );

    \I__1155\ : ClkMux
    port map (
            O => \N__5743\,
            I => \N__5595\
        );

    \I__1154\ : ClkMux
    port map (
            O => \N__5742\,
            I => \N__5595\
        );

    \I__1153\ : ClkMux
    port map (
            O => \N__5741\,
            I => \N__5595\
        );

    \I__1152\ : ClkMux
    port map (
            O => \N__5740\,
            I => \N__5595\
        );

    \I__1151\ : ClkMux
    port map (
            O => \N__5739\,
            I => \N__5595\
        );

    \I__1150\ : ClkMux
    port map (
            O => \N__5738\,
            I => \N__5595\
        );

    \I__1149\ : ClkMux
    port map (
            O => \N__5737\,
            I => \N__5595\
        );

    \I__1148\ : ClkMux
    port map (
            O => \N__5736\,
            I => \N__5595\
        );

    \I__1147\ : ClkMux
    port map (
            O => \N__5735\,
            I => \N__5595\
        );

    \I__1146\ : ClkMux
    port map (
            O => \N__5734\,
            I => \N__5595\
        );

    \I__1145\ : ClkMux
    port map (
            O => \N__5733\,
            I => \N__5595\
        );

    \I__1144\ : ClkMux
    port map (
            O => \N__5732\,
            I => \N__5595\
        );

    \I__1143\ : ClkMux
    port map (
            O => \N__5731\,
            I => \N__5595\
        );

    \I__1142\ : ClkMux
    port map (
            O => \N__5730\,
            I => \N__5595\
        );

    \I__1141\ : ClkMux
    port map (
            O => \N__5729\,
            I => \N__5595\
        );

    \I__1140\ : ClkMux
    port map (
            O => \N__5728\,
            I => \N__5595\
        );

    \I__1139\ : ClkMux
    port map (
            O => \N__5727\,
            I => \N__5595\
        );

    \I__1138\ : ClkMux
    port map (
            O => \N__5726\,
            I => \N__5595\
        );

    \I__1137\ : ClkMux
    port map (
            O => \N__5725\,
            I => \N__5595\
        );

    \I__1136\ : ClkMux
    port map (
            O => \N__5724\,
            I => \N__5595\
        );

    \I__1135\ : ClkMux
    port map (
            O => \N__5723\,
            I => \N__5595\
        );

    \I__1134\ : ClkMux
    port map (
            O => \N__5722\,
            I => \N__5595\
        );

    \I__1133\ : ClkMux
    port map (
            O => \N__5721\,
            I => \N__5595\
        );

    \I__1132\ : ClkMux
    port map (
            O => \N__5720\,
            I => \N__5595\
        );

    \I__1131\ : ClkMux
    port map (
            O => \N__5719\,
            I => \N__5595\
        );

    \I__1130\ : ClkMux
    port map (
            O => \N__5718\,
            I => \N__5595\
        );

    \I__1129\ : ClkMux
    port map (
            O => \N__5717\,
            I => \N__5595\
        );

    \I__1128\ : ClkMux
    port map (
            O => \N__5716\,
            I => \N__5595\
        );

    \I__1127\ : ClkMux
    port map (
            O => \N__5715\,
            I => \N__5595\
        );

    \I__1126\ : ClkMux
    port map (
            O => \N__5714\,
            I => \N__5595\
        );

    \I__1125\ : ClkMux
    port map (
            O => \N__5713\,
            I => \N__5595\
        );

    \I__1124\ : ClkMux
    port map (
            O => \N__5712\,
            I => \N__5595\
        );

    \I__1123\ : ClkMux
    port map (
            O => \N__5711\,
            I => \N__5595\
        );

    \I__1122\ : ClkMux
    port map (
            O => \N__5710\,
            I => \N__5595\
        );

    \I__1121\ : GlobalMux
    port map (
            O => \N__5595\,
            I => \N__5592\
        );

    \I__1120\ : gio2CtrlBuf
    port map (
            O => \N__5592\,
            I => \CLK_c_g\
        );

    \I__1119\ : CEMux
    port map (
            O => \N__5589\,
            I => \N__5496\
        );

    \I__1118\ : CEMux
    port map (
            O => \N__5588\,
            I => \N__5496\
        );

    \I__1117\ : CEMux
    port map (
            O => \N__5587\,
            I => \N__5496\
        );

    \I__1116\ : CEMux
    port map (
            O => \N__5586\,
            I => \N__5496\
        );

    \I__1115\ : CEMux
    port map (
            O => \N__5585\,
            I => \N__5496\
        );

    \I__1114\ : CEMux
    port map (
            O => \N__5584\,
            I => \N__5496\
        );

    \I__1113\ : CEMux
    port map (
            O => \N__5583\,
            I => \N__5496\
        );

    \I__1112\ : CEMux
    port map (
            O => \N__5582\,
            I => \N__5496\
        );

    \I__1111\ : CEMux
    port map (
            O => \N__5581\,
            I => \N__5496\
        );

    \I__1110\ : CEMux
    port map (
            O => \N__5580\,
            I => \N__5496\
        );

    \I__1109\ : CEMux
    port map (
            O => \N__5579\,
            I => \N__5496\
        );

    \I__1108\ : CEMux
    port map (
            O => \N__5578\,
            I => \N__5496\
        );

    \I__1107\ : CEMux
    port map (
            O => \N__5577\,
            I => \N__5496\
        );

    \I__1106\ : CEMux
    port map (
            O => \N__5576\,
            I => \N__5496\
        );

    \I__1105\ : CEMux
    port map (
            O => \N__5575\,
            I => \N__5496\
        );

    \I__1104\ : CEMux
    port map (
            O => \N__5574\,
            I => \N__5496\
        );

    \I__1103\ : CEMux
    port map (
            O => \N__5573\,
            I => \N__5496\
        );

    \I__1102\ : CEMux
    port map (
            O => \N__5572\,
            I => \N__5496\
        );

    \I__1101\ : CEMux
    port map (
            O => \N__5571\,
            I => \N__5496\
        );

    \I__1100\ : CEMux
    port map (
            O => \N__5570\,
            I => \N__5496\
        );

    \I__1099\ : CEMux
    port map (
            O => \N__5569\,
            I => \N__5496\
        );

    \I__1098\ : CEMux
    port map (
            O => \N__5568\,
            I => \N__5496\
        );

    \I__1097\ : CEMux
    port map (
            O => \N__5567\,
            I => \N__5496\
        );

    \I__1096\ : CEMux
    port map (
            O => \N__5566\,
            I => \N__5496\
        );

    \I__1095\ : CEMux
    port map (
            O => \N__5565\,
            I => \N__5496\
        );

    \I__1094\ : CEMux
    port map (
            O => \N__5564\,
            I => \N__5496\
        );

    \I__1093\ : CEMux
    port map (
            O => \N__5563\,
            I => \N__5496\
        );

    \I__1092\ : CEMux
    port map (
            O => \N__5562\,
            I => \N__5496\
        );

    \I__1091\ : CEMux
    port map (
            O => \N__5561\,
            I => \N__5496\
        );

    \I__1090\ : CEMux
    port map (
            O => \N__5560\,
            I => \N__5496\
        );

    \I__1089\ : CEMux
    port map (
            O => \N__5559\,
            I => \N__5496\
        );

    \I__1088\ : GlobalMux
    port map (
            O => \N__5496\,
            I => \N__5493\
        );

    \I__1087\ : gio2CtrlBuf
    port map (
            O => \N__5493\,
            I => \SEL_REG_i_g\
        );

    \I__1086\ : SRMux
    port map (
            O => \N__5490\,
            I => \N__5319\
        );

    \I__1085\ : SRMux
    port map (
            O => \N__5489\,
            I => \N__5319\
        );

    \I__1084\ : SRMux
    port map (
            O => \N__5488\,
            I => \N__5319\
        );

    \I__1083\ : SRMux
    port map (
            O => \N__5487\,
            I => \N__5319\
        );

    \I__1082\ : SRMux
    port map (
            O => \N__5486\,
            I => \N__5319\
        );

    \I__1081\ : SRMux
    port map (
            O => \N__5485\,
            I => \N__5319\
        );

    \I__1080\ : SRMux
    port map (
            O => \N__5484\,
            I => \N__5319\
        );

    \I__1079\ : SRMux
    port map (
            O => \N__5483\,
            I => \N__5319\
        );

    \I__1078\ : SRMux
    port map (
            O => \N__5482\,
            I => \N__5319\
        );

    \I__1077\ : SRMux
    port map (
            O => \N__5481\,
            I => \N__5319\
        );

    \I__1076\ : SRMux
    port map (
            O => \N__5480\,
            I => \N__5319\
        );

    \I__1075\ : SRMux
    port map (
            O => \N__5479\,
            I => \N__5319\
        );

    \I__1074\ : SRMux
    port map (
            O => \N__5478\,
            I => \N__5319\
        );

    \I__1073\ : SRMux
    port map (
            O => \N__5477\,
            I => \N__5319\
        );

    \I__1072\ : SRMux
    port map (
            O => \N__5476\,
            I => \N__5319\
        );

    \I__1071\ : SRMux
    port map (
            O => \N__5475\,
            I => \N__5319\
        );

    \I__1070\ : SRMux
    port map (
            O => \N__5474\,
            I => \N__5319\
        );

    \I__1069\ : SRMux
    port map (
            O => \N__5473\,
            I => \N__5319\
        );

    \I__1068\ : SRMux
    port map (
            O => \N__5472\,
            I => \N__5319\
        );

    \I__1067\ : SRMux
    port map (
            O => \N__5471\,
            I => \N__5319\
        );

    \I__1066\ : SRMux
    port map (
            O => \N__5470\,
            I => \N__5319\
        );

    \I__1065\ : SRMux
    port map (
            O => \N__5469\,
            I => \N__5319\
        );

    \I__1064\ : SRMux
    port map (
            O => \N__5468\,
            I => \N__5319\
        );

    \I__1063\ : SRMux
    port map (
            O => \N__5467\,
            I => \N__5319\
        );

    \I__1062\ : SRMux
    port map (
            O => \N__5466\,
            I => \N__5319\
        );

    \I__1061\ : SRMux
    port map (
            O => \N__5465\,
            I => \N__5319\
        );

    \I__1060\ : SRMux
    port map (
            O => \N__5464\,
            I => \N__5319\
        );

    \I__1059\ : SRMux
    port map (
            O => \N__5463\,
            I => \N__5319\
        );

    \I__1058\ : SRMux
    port map (
            O => \N__5462\,
            I => \N__5319\
        );

    \I__1057\ : SRMux
    port map (
            O => \N__5461\,
            I => \N__5319\
        );

    \I__1056\ : SRMux
    port map (
            O => \N__5460\,
            I => \N__5319\
        );

    \I__1055\ : SRMux
    port map (
            O => \N__5459\,
            I => \N__5319\
        );

    \I__1054\ : SRMux
    port map (
            O => \N__5458\,
            I => \N__5319\
        );

    \I__1053\ : SRMux
    port map (
            O => \N__5457\,
            I => \N__5319\
        );

    \I__1052\ : SRMux
    port map (
            O => \N__5456\,
            I => \N__5319\
        );

    \I__1051\ : SRMux
    port map (
            O => \N__5455\,
            I => \N__5319\
        );

    \I__1050\ : SRMux
    port map (
            O => \N__5454\,
            I => \N__5319\
        );

    \I__1049\ : SRMux
    port map (
            O => \N__5453\,
            I => \N__5319\
        );

    \I__1048\ : SRMux
    port map (
            O => \N__5452\,
            I => \N__5319\
        );

    \I__1047\ : SRMux
    port map (
            O => \N__5451\,
            I => \N__5319\
        );

    \I__1046\ : SRMux
    port map (
            O => \N__5450\,
            I => \N__5319\
        );

    \I__1045\ : SRMux
    port map (
            O => \N__5449\,
            I => \N__5319\
        );

    \I__1044\ : SRMux
    port map (
            O => \N__5448\,
            I => \N__5319\
        );

    \I__1043\ : SRMux
    port map (
            O => \N__5447\,
            I => \N__5319\
        );

    \I__1042\ : SRMux
    port map (
            O => \N__5446\,
            I => \N__5319\
        );

    \I__1041\ : SRMux
    port map (
            O => \N__5445\,
            I => \N__5319\
        );

    \I__1040\ : SRMux
    port map (
            O => \N__5444\,
            I => \N__5319\
        );

    \I__1039\ : SRMux
    port map (
            O => \N__5443\,
            I => \N__5319\
        );

    \I__1038\ : SRMux
    port map (
            O => \N__5442\,
            I => \N__5319\
        );

    \I__1037\ : SRMux
    port map (
            O => \N__5441\,
            I => \N__5319\
        );

    \I__1036\ : SRMux
    port map (
            O => \N__5440\,
            I => \N__5319\
        );

    \I__1035\ : SRMux
    port map (
            O => \N__5439\,
            I => \N__5319\
        );

    \I__1034\ : SRMux
    port map (
            O => \N__5438\,
            I => \N__5319\
        );

    \I__1033\ : SRMux
    port map (
            O => \N__5437\,
            I => \N__5319\
        );

    \I__1032\ : SRMux
    port map (
            O => \N__5436\,
            I => \N__5319\
        );

    \I__1031\ : SRMux
    port map (
            O => \N__5435\,
            I => \N__5319\
        );

    \I__1030\ : SRMux
    port map (
            O => \N__5434\,
            I => \N__5319\
        );

    \I__1029\ : GlobalMux
    port map (
            O => \N__5319\,
            I => \N__5316\
        );

    \I__1028\ : gio2CtrlBuf
    port map (
            O => \N__5316\,
            I => \RST_N_c_i_g\
        );

    \I__1027\ : InMux
    port map (
            O => \N__5313\,
            I => \N__5310\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__5310\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_57\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5307\,
            I => \N__5304\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__5304\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_58\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5301\,
            I => \N__5298\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__5298\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_61\
        );

    \I__1021\ : InMux
    port map (
            O => \N__5295\,
            I => \N__5292\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__5292\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_62\
        );

    \I__1019\ : InMux
    port map (
            O => \N__5289\,
            I => \N__5286\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5286\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_63\
        );

    \I__1017\ : InMux
    port map (
            O => \N__5283\,
            I => \N__5280\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__5280\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_64\
        );

    \I__1015\ : InMux
    port map (
            O => \N__5277\,
            I => \N__5274\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5274\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_65\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5271\,
            I => \N__5268\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5268\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_46\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5265\,
            I => \N__5262\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__5262\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_44\
        );

    \I__1009\ : InMux
    port map (
            O => \N__5259\,
            I => \N__5256\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5256\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_45\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5253\,
            I => \N__5250\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__5250\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_39\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5247\,
            I => \N__5244\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__5244\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_40\
        );

    \I__1003\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5238\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__5238\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_41\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5235\,
            I => \N__5232\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__5232\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_42\
        );

    \I__999\ : InMux
    port map (
            O => \N__5229\,
            I => \N__5226\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__5226\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_43\
        );

    \I__997\ : InMux
    port map (
            O => \N__5223\,
            I => \N__5220\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5220\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_59\
        );

    \I__995\ : InMux
    port map (
            O => \N__5217\,
            I => \N__5214\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5214\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_60\
        );

    \I__993\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5208\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__5208\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_72\
        );

    \I__991\ : InMux
    port map (
            O => \N__5205\,
            I => \N__5202\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__5202\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_35\
        );

    \I__989\ : InMux
    port map (
            O => \N__5199\,
            I => \N__5196\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__5196\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_36\
        );

    \I__987\ : InMux
    port map (
            O => \N__5193\,
            I => \N__5190\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__5190\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_37\
        );

    \I__985\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5184\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__5184\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_38\
        );

    \I__983\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5178\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5178\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_70\
        );

    \I__981\ : InMux
    port map (
            O => \N__5175\,
            I => \N__5172\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__5172\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_66\
        );

    \I__979\ : InMux
    port map (
            O => \N__5169\,
            I => \N__5166\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5166\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_67\
        );

    \I__977\ : InMux
    port map (
            O => \N__5163\,
            I => \N__5160\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__5160\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_68\
        );

    \I__975\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5154\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__5154\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_69\
        );

    \I__973\ : InMux
    port map (
            O => \N__5151\,
            I => \N__5148\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__5148\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_78\
        );

    \I__971\ : InMux
    port map (
            O => \N__5145\,
            I => \N__5142\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__5142\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_21\
        );

    \I__969\ : InMux
    port map (
            O => \N__5139\,
            I => \N__5136\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5136\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_22\
        );

    \I__967\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5130\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5130\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_19\
        );

    \I__965\ : InMux
    port map (
            O => \N__5127\,
            I => \N__5124\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__5124\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_20\
        );

    \I__963\ : InMux
    port map (
            O => \N__5121\,
            I => \N__5118\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__5118\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_75\
        );

    \I__961\ : InMux
    port map (
            O => \N__5115\,
            I => \N__5112\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__5112\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_76\
        );

    \I__959\ : InMux
    port map (
            O => \N__5109\,
            I => \N__5106\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__5106\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_77\
        );

    \I__957\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5100\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__5100\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_73\
        );

    \I__955\ : InMux
    port map (
            O => \N__5097\,
            I => \N__5094\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__5094\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_74\
        );

    \I__953\ : InMux
    port map (
            O => \N__5091\,
            I => \N__5088\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__5088\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_71\
        );

    \I__951\ : InMux
    port map (
            O => \N__5085\,
            I => \N__5082\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__5082\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_28\
        );

    \I__949\ : InMux
    port map (
            O => \N__5079\,
            I => \N__5076\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__5076\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_29\
        );

    \I__947\ : InMux
    port map (
            O => \N__5073\,
            I => \N__5070\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__5070\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_25\
        );

    \I__945\ : InMux
    port map (
            O => \N__5067\,
            I => \N__5064\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__5064\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_26\
        );

    \I__943\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5058\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__5058\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_34\
        );

    \I__941\ : InMux
    port map (
            O => \N__5055\,
            I => \N__5052\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__5052\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_23\
        );

    \I__939\ : InMux
    port map (
            O => \N__5049\,
            I => \N__5046\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5046\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_24\
        );

    \I__937\ : InMux
    port map (
            O => \N__5043\,
            I => \N__5040\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__5040\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_79\
        );

    \I__935\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5034\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5034\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_18\
        );

    \I__933\ : InMux
    port map (
            O => \N__5031\,
            I => \N__5028\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__5028\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_17\
        );

    \I__931\ : InMux
    port map (
            O => \N__5025\,
            I => \N__5022\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__5022\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_80\
        );

    \I__929\ : InMux
    port map (
            O => \N__5019\,
            I => \N__5016\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__5016\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_33\
        );

    \I__927\ : InMux
    port map (
            O => \N__5013\,
            I => \N__5010\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__5010\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_32\
        );

    \I__925\ : InMux
    port map (
            O => \N__5007\,
            I => \N__5004\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5004\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_27\
        );

    \I__923\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4998\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__4998\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_30\
        );

    \I__921\ : InMux
    port map (
            O => \N__4995\,
            I => \N__4992\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4992\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_31\
        );

    \I__919\ : InMux
    port map (
            O => \N__4989\,
            I => \N__4986\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4986\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_15\
        );

    \I__917\ : InMux
    port map (
            O => \N__4983\,
            I => \N__4980\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4980\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_86\
        );

    \I__915\ : InMux
    port map (
            O => \N__4977\,
            I => \N__4974\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4974\,
            I => \N__4971\
        );

    \I__913\ : Span4Mux_v
    port map (
            O => \N__4971\,
            I => \N__4968\
        );

    \I__912\ : Span4Mux_h
    port map (
            O => \N__4968\,
            I => \N__4965\
        );

    \I__911\ : Odrv4
    port map (
            O => \N__4965\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_87\
        );

    \I__910\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4959\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__4959\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_85\
        );

    \I__908\ : InMux
    port map (
            O => \N__4956\,
            I => \N__4953\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__4953\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_84\
        );

    \I__906\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4947\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__4947\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_83\
        );

    \I__904\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4941\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4941\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_16\
        );

    \I__902\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4935\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4935\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_82\
        );

    \I__900\ : InMux
    port map (
            O => \N__4932\,
            I => \N__4929\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__4929\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_81\
        );

    \I__898\ : InMux
    port map (
            O => \N__4926\,
            I => \N__4923\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__4923\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_6\
        );

    \I__896\ : InMux
    port map (
            O => \N__4920\,
            I => \N__4917\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4917\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_7\
        );

    \I__894\ : InMux
    port map (
            O => \N__4914\,
            I => \N__4911\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4911\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_10\
        );

    \I__892\ : InMux
    port map (
            O => \N__4908\,
            I => \N__4905\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__4905\,
            I => \N__4902\
        );

    \I__890\ : Odrv4
    port map (
            O => \N__4902\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_8\
        );

    \I__889\ : InMux
    port map (
            O => \N__4899\,
            I => \N__4896\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__4896\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_9\
        );

    \I__887\ : InMux
    port map (
            O => \N__4893\,
            I => \N__4890\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__4890\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_11\
        );

    \I__885\ : InMux
    port map (
            O => \N__4887\,
            I => \N__4884\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4884\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_12\
        );

    \I__883\ : InMux
    port map (
            O => \N__4881\,
            I => \N__4878\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4878\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_13\
        );

    \I__881\ : InMux
    port map (
            O => \N__4875\,
            I => \N__4872\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4872\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_14\
        );

    \I__879\ : InMux
    port map (
            O => \N__4869\,
            I => \N__4866\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__4866\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_12\
        );

    \I__877\ : InMux
    port map (
            O => \N__4863\,
            I => \N__4860\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4860\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_15\
        );

    \I__875\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4854\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__4854\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_13\
        );

    \I__873\ : InMux
    port map (
            O => \N__4851\,
            I => \N__4848\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4848\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_14\
        );

    \I__871\ : InMux
    port map (
            O => \N__4845\,
            I => \N__4842\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4842\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_7\
        );

    \I__869\ : InMux
    port map (
            O => \N__4839\,
            I => \N__4836\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4836\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_8\
        );

    \I__867\ : InMux
    port map (
            O => \N__4833\,
            I => \N__4830\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4830\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_9\
        );

    \I__865\ : InMux
    port map (
            O => \N__4827\,
            I => \N__4824\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4824\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_10\
        );

    \I__863\ : InMux
    port map (
            O => \N__4821\,
            I => \N__4818\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4818\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_11\
        );

    \I__861\ : CEMux
    port map (
            O => \N__4815\,
            I => \N__4811\
        );

    \I__860\ : CEMux
    port map (
            O => \N__4814\,
            I => \N__4807\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4811\,
            I => \N__4802\
        );

    \I__858\ : CEMux
    port map (
            O => \N__4810\,
            I => \N__4799\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4807\,
            I => \N__4796\
        );

    \I__856\ : CEMux
    port map (
            O => \N__4806\,
            I => \N__4793\
        );

    \I__855\ : InMux
    port map (
            O => \N__4805\,
            I => \N__4789\
        );

    \I__854\ : Span4Mux_v
    port map (
            O => \N__4802\,
            I => \N__4786\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4799\,
            I => \N__4783\
        );

    \I__852\ : Span4Mux_v
    port map (
            O => \N__4796\,
            I => \N__4780\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__4793\,
            I => \N__4777\
        );

    \I__850\ : InMux
    port map (
            O => \N__4792\,
            I => \N__4774\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__4789\,
            I => \SEL_REG\
        );

    \I__848\ : Odrv4
    port map (
            O => \N__4786\,
            I => \SEL_REG\
        );

    \I__847\ : Odrv4
    port map (
            O => \N__4783\,
            I => \SEL_REG\
        );

    \I__846\ : Odrv4
    port map (
            O => \N__4780\,
            I => \SEL_REG\
        );

    \I__845\ : Odrv12
    port map (
            O => \N__4777\,
            I => \SEL_REG\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__4774\,
            I => \SEL_REG\
        );

    \I__843\ : InMux
    port map (
            O => \N__4761\,
            I => \N__4758\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4758\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_4\
        );

    \I__841\ : InMux
    port map (
            O => \N__4755\,
            I => \N__4752\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4752\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_5\
        );

    \I__839\ : InMux
    port map (
            O => \N__4749\,
            I => \N__4741\
        );

    \I__838\ : InMux
    port map (
            O => \N__4748\,
            I => \N__4734\
        );

    \I__837\ : InMux
    port map (
            O => \N__4747\,
            I => \N__4734\
        );

    \I__836\ : InMux
    port map (
            O => \N__4746\,
            I => \N__4734\
        );

    \I__835\ : InMux
    port map (
            O => \N__4745\,
            I => \N__4729\
        );

    \I__834\ : InMux
    port map (
            O => \N__4744\,
            I => \N__4729\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4741\,
            I => \N__4711\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4734\,
            I => \N__4711\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4729\,
            I => \N__4711\
        );

    \I__830\ : InMux
    port map (
            O => \N__4728\,
            I => \N__4692\
        );

    \I__829\ : InMux
    port map (
            O => \N__4727\,
            I => \N__4692\
        );

    \I__828\ : InMux
    port map (
            O => \N__4726\,
            I => \N__4692\
        );

    \I__827\ : InMux
    port map (
            O => \N__4725\,
            I => \N__4692\
        );

    \I__826\ : InMux
    port map (
            O => \N__4724\,
            I => \N__4677\
        );

    \I__825\ : InMux
    port map (
            O => \N__4723\,
            I => \N__4677\
        );

    \I__824\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4677\
        );

    \I__823\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4677\
        );

    \I__822\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4677\
        );

    \I__821\ : InMux
    port map (
            O => \N__4719\,
            I => \N__4677\
        );

    \I__820\ : InMux
    port map (
            O => \N__4718\,
            I => \N__4677\
        );

    \I__819\ : Span4Mux_h
    port map (
            O => \N__4711\,
            I => \N__4674\
        );

    \I__818\ : InMux
    port map (
            O => \N__4710\,
            I => \N__4671\
        );

    \I__817\ : InMux
    port map (
            O => \N__4709\,
            I => \N__4658\
        );

    \I__816\ : InMux
    port map (
            O => \N__4708\,
            I => \N__4658\
        );

    \I__815\ : InMux
    port map (
            O => \N__4707\,
            I => \N__4658\
        );

    \I__814\ : InMux
    port map (
            O => \N__4706\,
            I => \N__4658\
        );

    \I__813\ : InMux
    port map (
            O => \N__4705\,
            I => \N__4658\
        );

    \I__812\ : InMux
    port map (
            O => \N__4704\,
            I => \N__4658\
        );

    \I__811\ : InMux
    port map (
            O => \N__4703\,
            I => \N__4651\
        );

    \I__810\ : InMux
    port map (
            O => \N__4702\,
            I => \N__4651\
        );

    \I__809\ : InMux
    port map (
            O => \N__4701\,
            I => \N__4651\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4692\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_0\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__4677\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_0\
        );

    \I__806\ : Odrv4
    port map (
            O => \N__4674\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_0\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__4671\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_0\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__4658\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_0\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__4651\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_0\
        );

    \I__802\ : IoInMux
    port map (
            O => \N__4638\,
            I => \N__4635\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__4635\,
            I => \N__4632\
        );

    \I__800\ : IoSpan4Mux
    port map (
            O => \N__4632\,
            I => \N__4629\
        );

    \I__799\ : Span4Mux_s0_v
    port map (
            O => \N__4629\,
            I => \N__4626\
        );

    \I__798\ : Sp12to4
    port map (
            O => \N__4626\,
            I => \N__4623\
        );

    \I__797\ : Span12Mux_s11_v
    port map (
            O => \N__4623\,
            I => \N__4620\
        );

    \I__796\ : Odrv12
    port map (
            O => \N__4620\,
            I => \fsm_ctrl_inst1.SEL_REG_i\
        );

    \I__795\ : InMux
    port map (
            O => \N__4617\,
            I => \N__4614\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__4614\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_4\
        );

    \I__793\ : InMux
    port map (
            O => \N__4611\,
            I => \N__4608\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__4608\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_5\
        );

    \I__791\ : InMux
    port map (
            O => \N__4605\,
            I => \N__4602\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4602\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_6\
        );

    \I__789\ : InMux
    port map (
            O => \N__4599\,
            I => \N__4596\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__4596\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_0\
        );

    \I__787\ : InMux
    port map (
            O => \N__4593\,
            I => \N__4590\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__4590\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_1\
        );

    \I__785\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4584\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__4584\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_2\
        );

    \I__783\ : InMux
    port map (
            O => \N__4581\,
            I => \N__4578\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__4578\,
            I => \config_register_latched_dec_inst1.STATSRZ0Z_3\
        );

    \I__781\ : InMux
    port map (
            O => \N__4575\,
            I => \N__4572\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__4572\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_0\
        );

    \I__779\ : InMux
    port map (
            O => \N__4569\,
            I => \N__4566\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__4566\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_2\
        );

    \I__777\ : InMux
    port map (
            O => \N__4563\,
            I => \N__4560\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__4560\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_3\
        );

    \I__775\ : InMux
    port map (
            O => \N__4557\,
            I => \N__4554\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4554\,
            I => \N__4550\
        );

    \I__773\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4547\
        );

    \I__772\ : Odrv4
    port map (
            O => \N__4550\,
            I => \MOSI\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__4547\,
            I => \MOSI\
        );

    \I__770\ : IoInMux
    port map (
            O => \N__4542\,
            I => \N__4539\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__4539\,
            I => \N__4536\
        );

    \I__768\ : IoSpan4Mux
    port map (
            O => \N__4536\,
            I => \N__4533\
        );

    \I__767\ : Sp12to4
    port map (
            O => \N__4533\,
            I => \N__4530\
        );

    \I__766\ : Span12Mux_s7_v
    port map (
            O => \N__4530\,
            I => \N__4527\
        );

    \I__765\ : Span12Mux_v
    port map (
            O => \N__4527\,
            I => \N__4524\
        );

    \I__764\ : Odrv12
    port map (
            O => \N__4524\,
            I => \SDO_signal_out_c\
        );

    \I__763\ : CascadeMux
    port map (
            O => \N__4521\,
            I => \fsm_ctrl_inst1.counter_din_RNO_0Z0Z_3_cascade_\
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__4518\,
            I => \N__4514\
        );

    \I__761\ : InMux
    port map (
            O => \N__4517\,
            I => \N__4509\
        );

    \I__760\ : InMux
    port map (
            O => \N__4514\,
            I => \N__4509\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__4509\,
            I => \fsm_ctrl_inst1.counter_dinZ0Z_3\
        );

    \I__758\ : InMux
    port map (
            O => \N__4506\,
            I => \N__4500\
        );

    \I__757\ : InMux
    port map (
            O => \N__4505\,
            I => \N__4500\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__4500\,
            I => \N__4497\
        );

    \I__755\ : Span4Mux_v
    port map (
            O => \N__4497\,
            I => \N__4493\
        );

    \I__754\ : InMux
    port map (
            O => \N__4496\,
            I => \N__4490\
        );

    \I__753\ : Odrv4
    port map (
            O => \N__4493\,
            I => \fsm_ctrl_inst1.counter_din_RNI6L3H1Z0Z_3\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__4490\,
            I => \fsm_ctrl_inst1.counter_din_RNI6L3H1Z0Z_3\
        );

    \I__751\ : CascadeMux
    port map (
            O => \N__4485\,
            I => \N__4481\
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__4484\,
            I => \N__4478\
        );

    \I__749\ : InMux
    port map (
            O => \N__4481\,
            I => \N__4470\
        );

    \I__748\ : InMux
    port map (
            O => \N__4478\,
            I => \N__4470\
        );

    \I__747\ : InMux
    port map (
            O => \N__4477\,
            I => \N__4470\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4470\,
            I => \fsm_ctrl_inst1.counter_dinZ0Z_2\
        );

    \I__745\ : CascadeMux
    port map (
            O => \N__4467\,
            I => \N__4462\
        );

    \I__744\ : InMux
    port map (
            O => \N__4466\,
            I => \N__4457\
        );

    \I__743\ : InMux
    port map (
            O => \N__4465\,
            I => \N__4448\
        );

    \I__742\ : InMux
    port map (
            O => \N__4462\,
            I => \N__4448\
        );

    \I__741\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4448\
        );

    \I__740\ : InMux
    port map (
            O => \N__4460\,
            I => \N__4448\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__4457\,
            I => \fsm_ctrl_inst1.counter_dinZ0Z_0\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4448\,
            I => \fsm_ctrl_inst1.counter_dinZ0Z_0\
        );

    \I__737\ : InMux
    port map (
            O => \N__4443\,
            I => \N__4431\
        );

    \I__736\ : InMux
    port map (
            O => \N__4442\,
            I => \N__4431\
        );

    \I__735\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4431\
        );

    \I__734\ : InMux
    port map (
            O => \N__4440\,
            I => \N__4431\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4431\,
            I => \fsm_ctrl_inst1.counter_dinZ0Z_1\
        );

    \I__732\ : InMux
    port map (
            O => \N__4428\,
            I => \N__4425\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4425\,
            I => \N__4422\
        );

    \I__730\ : Odrv12
    port map (
            O => \N__4422\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_83\
        );

    \I__729\ : InMux
    port map (
            O => \N__4419\,
            I => \N__4416\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__4416\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_84\
        );

    \I__727\ : InMux
    port map (
            O => \N__4413\,
            I => \N__4410\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__4410\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_85\
        );

    \I__725\ : InMux
    port map (
            O => \N__4407\,
            I => \N__4404\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__4404\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_86\
        );

    \I__723\ : CEMux
    port map (
            O => \N__4401\,
            I => \N__4359\
        );

    \I__722\ : CEMux
    port map (
            O => \N__4400\,
            I => \N__4359\
        );

    \I__721\ : CEMux
    port map (
            O => \N__4399\,
            I => \N__4359\
        );

    \I__720\ : CEMux
    port map (
            O => \N__4398\,
            I => \N__4359\
        );

    \I__719\ : CEMux
    port map (
            O => \N__4397\,
            I => \N__4359\
        );

    \I__718\ : CEMux
    port map (
            O => \N__4396\,
            I => \N__4359\
        );

    \I__717\ : CEMux
    port map (
            O => \N__4395\,
            I => \N__4359\
        );

    \I__716\ : CEMux
    port map (
            O => \N__4394\,
            I => \N__4359\
        );

    \I__715\ : CEMux
    port map (
            O => \N__4393\,
            I => \N__4359\
        );

    \I__714\ : CEMux
    port map (
            O => \N__4392\,
            I => \N__4359\
        );

    \I__713\ : CEMux
    port map (
            O => \N__4391\,
            I => \N__4359\
        );

    \I__712\ : CEMux
    port map (
            O => \N__4390\,
            I => \N__4359\
        );

    \I__711\ : CEMux
    port map (
            O => \N__4389\,
            I => \N__4359\
        );

    \I__710\ : CEMux
    port map (
            O => \N__4388\,
            I => \N__4359\
        );

    \I__709\ : GlobalMux
    port map (
            O => \N__4359\,
            I => \N__4356\
        );

    \I__708\ : gio2CtrlBuf
    port map (
            O => \N__4356\,
            I => \fsm_ctrl_inst1.current_state_i_g_0\
        );

    \I__707\ : InMux
    port map (
            O => \N__4353\,
            I => \N__4350\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4350\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_15\
        );

    \I__705\ : CascadeMux
    port map (
            O => \N__4347\,
            I => \N__4344\
        );

    \I__704\ : InMux
    port map (
            O => \N__4344\,
            I => \N__4341\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__4341\,
            I => \N__4338\
        );

    \I__702\ : Odrv4
    port map (
            O => \N__4338\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_87\
        );

    \I__701\ : InMux
    port map (
            O => \N__4335\,
            I => \N__4308\
        );

    \I__700\ : InMux
    port map (
            O => \N__4334\,
            I => \N__4295\
        );

    \I__699\ : InMux
    port map (
            O => \N__4333\,
            I => \N__4295\
        );

    \I__698\ : InMux
    port map (
            O => \N__4332\,
            I => \N__4295\
        );

    \I__697\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4295\
        );

    \I__696\ : InMux
    port map (
            O => \N__4330\,
            I => \N__4295\
        );

    \I__695\ : InMux
    port map (
            O => \N__4329\,
            I => \N__4295\
        );

    \I__694\ : InMux
    port map (
            O => \N__4328\,
            I => \N__4290\
        );

    \I__693\ : InMux
    port map (
            O => \N__4327\,
            I => \N__4290\
        );

    \I__692\ : InMux
    port map (
            O => \N__4326\,
            I => \N__4271\
        );

    \I__691\ : InMux
    port map (
            O => \N__4325\,
            I => \N__4271\
        );

    \I__690\ : InMux
    port map (
            O => \N__4324\,
            I => \N__4271\
        );

    \I__689\ : InMux
    port map (
            O => \N__4323\,
            I => \N__4271\
        );

    \I__688\ : InMux
    port map (
            O => \N__4322\,
            I => \N__4271\
        );

    \I__687\ : InMux
    port map (
            O => \N__4321\,
            I => \N__4229\
        );

    \I__686\ : InMux
    port map (
            O => \N__4320\,
            I => \N__4229\
        );

    \I__685\ : InMux
    port map (
            O => \N__4319\,
            I => \N__4229\
        );

    \I__684\ : InMux
    port map (
            O => \N__4318\,
            I => \N__4229\
        );

    \I__683\ : InMux
    port map (
            O => \N__4317\,
            I => \N__4222\
        );

    \I__682\ : InMux
    port map (
            O => \N__4316\,
            I => \N__4222\
        );

    \I__681\ : InMux
    port map (
            O => \N__4315\,
            I => \N__4222\
        );

    \I__680\ : InMux
    port map (
            O => \N__4314\,
            I => \N__4197\
        );

    \I__679\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4197\
        );

    \I__678\ : InMux
    port map (
            O => \N__4312\,
            I => \N__4197\
        );

    \I__677\ : InMux
    port map (
            O => \N__4311\,
            I => \N__4197\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__4308\,
            I => \N__4194\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__4295\,
            I => \N__4191\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__4290\,
            I => \N__4188\
        );

    \I__673\ : InMux
    port map (
            O => \N__4289\,
            I => \N__4171\
        );

    \I__672\ : InMux
    port map (
            O => \N__4288\,
            I => \N__4171\
        );

    \I__671\ : InMux
    port map (
            O => \N__4287\,
            I => \N__4171\
        );

    \I__670\ : InMux
    port map (
            O => \N__4286\,
            I => \N__4171\
        );

    \I__669\ : InMux
    port map (
            O => \N__4285\,
            I => \N__4171\
        );

    \I__668\ : InMux
    port map (
            O => \N__4284\,
            I => \N__4171\
        );

    \I__667\ : InMux
    port map (
            O => \N__4283\,
            I => \N__4171\
        );

    \I__666\ : InMux
    port map (
            O => \N__4282\,
            I => \N__4171\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__4271\,
            I => \N__4168\
        );

    \I__664\ : InMux
    port map (
            O => \N__4270\,
            I => \N__4151\
        );

    \I__663\ : InMux
    port map (
            O => \N__4269\,
            I => \N__4151\
        );

    \I__662\ : InMux
    port map (
            O => \N__4268\,
            I => \N__4151\
        );

    \I__661\ : InMux
    port map (
            O => \N__4267\,
            I => \N__4151\
        );

    \I__660\ : InMux
    port map (
            O => \N__4266\,
            I => \N__4151\
        );

    \I__659\ : InMux
    port map (
            O => \N__4265\,
            I => \N__4151\
        );

    \I__658\ : InMux
    port map (
            O => \N__4264\,
            I => \N__4151\
        );

    \I__657\ : InMux
    port map (
            O => \N__4263\,
            I => \N__4151\
        );

    \I__656\ : InMux
    port map (
            O => \N__4262\,
            I => \N__4134\
        );

    \I__655\ : InMux
    port map (
            O => \N__4261\,
            I => \N__4134\
        );

    \I__654\ : InMux
    port map (
            O => \N__4260\,
            I => \N__4134\
        );

    \I__653\ : InMux
    port map (
            O => \N__4259\,
            I => \N__4134\
        );

    \I__652\ : InMux
    port map (
            O => \N__4258\,
            I => \N__4134\
        );

    \I__651\ : InMux
    port map (
            O => \N__4257\,
            I => \N__4134\
        );

    \I__650\ : InMux
    port map (
            O => \N__4256\,
            I => \N__4134\
        );

    \I__649\ : InMux
    port map (
            O => \N__4255\,
            I => \N__4134\
        );

    \I__648\ : InMux
    port map (
            O => \N__4254\,
            I => \N__4117\
        );

    \I__647\ : InMux
    port map (
            O => \N__4253\,
            I => \N__4117\
        );

    \I__646\ : InMux
    port map (
            O => \N__4252\,
            I => \N__4117\
        );

    \I__645\ : InMux
    port map (
            O => \N__4251\,
            I => \N__4117\
        );

    \I__644\ : InMux
    port map (
            O => \N__4250\,
            I => \N__4117\
        );

    \I__643\ : InMux
    port map (
            O => \N__4249\,
            I => \N__4117\
        );

    \I__642\ : InMux
    port map (
            O => \N__4248\,
            I => \N__4117\
        );

    \I__641\ : InMux
    port map (
            O => \N__4247\,
            I => \N__4117\
        );

    \I__640\ : InMux
    port map (
            O => \N__4246\,
            I => \N__4100\
        );

    \I__639\ : InMux
    port map (
            O => \N__4245\,
            I => \N__4100\
        );

    \I__638\ : InMux
    port map (
            O => \N__4244\,
            I => \N__4100\
        );

    \I__637\ : InMux
    port map (
            O => \N__4243\,
            I => \N__4100\
        );

    \I__636\ : InMux
    port map (
            O => \N__4242\,
            I => \N__4100\
        );

    \I__635\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4100\
        );

    \I__634\ : InMux
    port map (
            O => \N__4240\,
            I => \N__4100\
        );

    \I__633\ : InMux
    port map (
            O => \N__4239\,
            I => \N__4100\
        );

    \I__632\ : CascadeMux
    port map (
            O => \N__4238\,
            I => \N__4088\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__4229\,
            I => \N__4081\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4222\,
            I => \N__4078\
        );

    \I__629\ : InMux
    port map (
            O => \N__4221\,
            I => \N__4061\
        );

    \I__628\ : InMux
    port map (
            O => \N__4220\,
            I => \N__4061\
        );

    \I__627\ : InMux
    port map (
            O => \N__4219\,
            I => \N__4061\
        );

    \I__626\ : InMux
    port map (
            O => \N__4218\,
            I => \N__4061\
        );

    \I__625\ : InMux
    port map (
            O => \N__4217\,
            I => \N__4061\
        );

    \I__624\ : InMux
    port map (
            O => \N__4216\,
            I => \N__4061\
        );

    \I__623\ : InMux
    port map (
            O => \N__4215\,
            I => \N__4061\
        );

    \I__622\ : InMux
    port map (
            O => \N__4214\,
            I => \N__4061\
        );

    \I__621\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4044\
        );

    \I__620\ : InMux
    port map (
            O => \N__4212\,
            I => \N__4044\
        );

    \I__619\ : InMux
    port map (
            O => \N__4211\,
            I => \N__4044\
        );

    \I__618\ : InMux
    port map (
            O => \N__4210\,
            I => \N__4044\
        );

    \I__617\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4044\
        );

    \I__616\ : InMux
    port map (
            O => \N__4208\,
            I => \N__4044\
        );

    \I__615\ : InMux
    port map (
            O => \N__4207\,
            I => \N__4044\
        );

    \I__614\ : InMux
    port map (
            O => \N__4206\,
            I => \N__4044\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__4197\,
            I => \N__4041\
        );

    \I__612\ : Span4Mux_v
    port map (
            O => \N__4194\,
            I => \N__4032\
        );

    \I__611\ : Span4Mux_v
    port map (
            O => \N__4191\,
            I => \N__4032\
        );

    \I__610\ : Span4Mux_v
    port map (
            O => \N__4188\,
            I => \N__4032\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__4171\,
            I => \N__4032\
        );

    \I__608\ : Span4Mux_s2_h
    port map (
            O => \N__4168\,
            I => \N__4025\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__4151\,
            I => \N__4025\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__4134\,
            I => \N__4025\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__4117\,
            I => \N__4020\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__4100\,
            I => \N__4020\
        );

    \I__603\ : InMux
    port map (
            O => \N__4099\,
            I => \N__4003\
        );

    \I__602\ : InMux
    port map (
            O => \N__4098\,
            I => \N__4003\
        );

    \I__601\ : InMux
    port map (
            O => \N__4097\,
            I => \N__4003\
        );

    \I__600\ : InMux
    port map (
            O => \N__4096\,
            I => \N__4003\
        );

    \I__599\ : InMux
    port map (
            O => \N__4095\,
            I => \N__4003\
        );

    \I__598\ : InMux
    port map (
            O => \N__4094\,
            I => \N__4003\
        );

    \I__597\ : InMux
    port map (
            O => \N__4093\,
            I => \N__4003\
        );

    \I__596\ : InMux
    port map (
            O => \N__4092\,
            I => \N__4003\
        );

    \I__595\ : InMux
    port map (
            O => \N__4091\,
            I => \N__3996\
        );

    \I__594\ : InMux
    port map (
            O => \N__4088\,
            I => \N__3996\
        );

    \I__593\ : InMux
    port map (
            O => \N__4087\,
            I => \N__3996\
        );

    \I__592\ : InMux
    port map (
            O => \N__4086\,
            I => \N__3993\
        );

    \I__591\ : InMux
    port map (
            O => \N__4085\,
            I => \N__3988\
        );

    \I__590\ : InMux
    port map (
            O => \N__4084\,
            I => \N__3988\
        );

    \I__589\ : Odrv4
    port map (
            O => \N__4081\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__588\ : Odrv4
    port map (
            O => \N__4078\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4061\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4044\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__585\ : Odrv4
    port map (
            O => \N__4041\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__584\ : Odrv4
    port map (
            O => \N__4032\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__583\ : Odrv4
    port map (
            O => \N__4025\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__582\ : Odrv4
    port map (
            O => \N__4020\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__4003\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3996\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__3993\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3988\,
            I => \fsm_ctrl_inst1.current_stateZ0Z_1\
        );

    \I__577\ : InMux
    port map (
            O => \N__3963\,
            I => \N__3960\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3960\,
            I => \config_register_latched_dec_inst1.DYNSRZ0Z_1\
        );

    \I__575\ : InMux
    port map (
            O => \N__3957\,
            I => \N__3954\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__3954\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_12\
        );

    \I__573\ : InMux
    port map (
            O => \N__3951\,
            I => \N__3948\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3948\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_13\
        );

    \I__571\ : InMux
    port map (
            O => \N__3945\,
            I => \N__3942\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3942\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_14\
        );

    \I__569\ : InMux
    port map (
            O => \N__3939\,
            I => \N__3936\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3936\,
            I => \N__3933\
        );

    \I__567\ : Odrv4
    port map (
            O => \N__3933\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_8\
        );

    \I__566\ : InMux
    port map (
            O => \N__3930\,
            I => \N__3927\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__3927\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_9\
        );

    \I__564\ : CEMux
    port map (
            O => \N__3924\,
            I => \N__3921\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3921\,
            I => \N__3916\
        );

    \I__562\ : CEMux
    port map (
            O => \N__3920\,
            I => \N__3913\
        );

    \I__561\ : CEMux
    port map (
            O => \N__3919\,
            I => \N__3910\
        );

    \I__560\ : Odrv12
    port map (
            O => \N__3916\,
            I => \fsm_ctrl_inst1.current_state_i_1\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3913\,
            I => \fsm_ctrl_inst1.current_state_i_1\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__3910\,
            I => \fsm_ctrl_inst1.current_state_i_1\
        );

    \I__557\ : InMux
    port map (
            O => \N__3903\,
            I => \N__3900\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__3900\,
            I => \N__3897\
        );

    \I__555\ : Odrv12
    port map (
            O => \N__3897\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_46\
        );

    \I__554\ : InMux
    port map (
            O => \N__3894\,
            I => \N__3891\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3891\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_47\
        );

    \I__552\ : InMux
    port map (
            O => \N__3888\,
            I => \N__3885\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3885\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_53\
        );

    \I__550\ : InMux
    port map (
            O => \N__3882\,
            I => \N__3879\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3879\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_52\
        );

    \I__548\ : InMux
    port map (
            O => \N__3876\,
            I => \N__3873\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3873\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_50\
        );

    \I__546\ : InMux
    port map (
            O => \N__3870\,
            I => \N__3867\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3867\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_51\
        );

    \I__544\ : InMux
    port map (
            O => \N__3864\,
            I => \N__3861\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3861\,
            I => \CONSTANT_ONE_NET\
        );

    \I__542\ : InMux
    port map (
            O => \N__3858\,
            I => \N__3855\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3855\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_4\
        );

    \I__540\ : InMux
    port map (
            O => \N__3852\,
            I => \N__3849\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3849\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_5\
        );

    \I__538\ : InMux
    port map (
            O => \N__3846\,
            I => \N__3843\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3843\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_6\
        );

    \I__536\ : InMux
    port map (
            O => \N__3840\,
            I => \N__3837\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3837\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_7\
        );

    \I__534\ : CEMux
    port map (
            O => \N__3834\,
            I => \N__3831\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3831\,
            I => \N__3823\
        );

    \I__532\ : InMux
    port map (
            O => \N__3830\,
            I => \N__3818\
        );

    \I__531\ : InMux
    port map (
            O => \N__3829\,
            I => \N__3818\
        );

    \I__530\ : InMux
    port map (
            O => \N__3828\,
            I => \N__3811\
        );

    \I__529\ : InMux
    port map (
            O => \N__3827\,
            I => \N__3811\
        );

    \I__528\ : InMux
    port map (
            O => \N__3826\,
            I => \N__3811\
        );

    \I__527\ : Span4Mux_s3_h
    port map (
            O => \N__3823\,
            I => \N__3808\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3818\,
            I => \fsm_ctrl_inst1.counter_state_0_i\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3811\,
            I => \fsm_ctrl_inst1.counter_state_0_i\
        );

    \I__524\ : Odrv4
    port map (
            O => \N__3808\,
            I => \fsm_ctrl_inst1.counter_state_0_i\
        );

    \I__523\ : InMux
    port map (
            O => \N__3801\,
            I => \N__3797\
        );

    \I__522\ : InMux
    port map (
            O => \N__3800\,
            I => \N__3794\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3797\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_3\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3794\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_3\
        );

    \I__519\ : InMux
    port map (
            O => \N__3789\,
            I => \N__3785\
        );

    \I__518\ : InMux
    port map (
            O => \N__3788\,
            I => \N__3782\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3785\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_2\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3782\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_2\
        );

    \I__515\ : InMux
    port map (
            O => \N__3777\,
            I => \N__3773\
        );

    \I__514\ : InMux
    port map (
            O => \N__3776\,
            I => \N__3770\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3773\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_4\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3770\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_4\
        );

    \I__511\ : InMux
    port map (
            O => \N__3765\,
            I => \N__3759\
        );

    \I__510\ : InMux
    port map (
            O => \N__3764\,
            I => \N__3759\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3759\,
            I => \fsm_ctrl_inst1.N_127_1\
        );

    \I__508\ : InMux
    port map (
            O => \N__3756\,
            I => \N__3753\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3753\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_10\
        );

    \I__506\ : InMux
    port map (
            O => \N__3750\,
            I => \N__3747\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3747\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_11\
        );

    \I__504\ : InMux
    port map (
            O => \N__3744\,
            I => \N__3741\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3741\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_44\
        );

    \I__502\ : InMux
    port map (
            O => \N__3738\,
            I => \N__3733\
        );

    \I__501\ : InMux
    port map (
            O => \N__3737\,
            I => \N__3730\
        );

    \I__500\ : InMux
    port map (
            O => \N__3736\,
            I => \N__3727\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3733\,
            I => \N__3724\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3730\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_4\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3727\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_4\
        );

    \I__496\ : Odrv4
    port map (
            O => \N__3724\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_4\
        );

    \I__495\ : InMux
    port map (
            O => \N__3717\,
            I => \N__3712\
        );

    \I__494\ : InMux
    port map (
            O => \N__3716\,
            I => \N__3709\
        );

    \I__493\ : InMux
    port map (
            O => \N__3715\,
            I => \N__3706\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3712\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_3\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3709\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_3\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3706\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_3\
        );

    \I__489\ : CascadeMux
    port map (
            O => \N__3699\,
            I => \N__3696\
        );

    \I__488\ : InMux
    port map (
            O => \N__3696\,
            I => \N__3691\
        );

    \I__487\ : InMux
    port map (
            O => \N__3695\,
            I => \N__3688\
        );

    \I__486\ : InMux
    port map (
            O => \N__3694\,
            I => \N__3685\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3691\,
            I => \N__3682\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3688\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_5\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__3685\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_5\
        );

    \I__482\ : Odrv4
    port map (
            O => \N__3682\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_5\
        );

    \I__481\ : InMux
    port map (
            O => \N__3675\,
            I => \N__3670\
        );

    \I__480\ : InMux
    port map (
            O => \N__3674\,
            I => \N__3667\
        );

    \I__479\ : InMux
    port map (
            O => \N__3673\,
            I => \N__3664\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__3670\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_6\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3667\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_6\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3664\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_6\
        );

    \I__475\ : CascadeMux
    port map (
            O => \N__3657\,
            I => \fsm_ctrl_inst1.counter_stat_RNIML9Z0Z_6_cascade_\
        );

    \I__474\ : InMux
    port map (
            O => \N__3654\,
            I => \N__3642\
        );

    \I__473\ : InMux
    port map (
            O => \N__3653\,
            I => \N__3642\
        );

    \I__472\ : InMux
    port map (
            O => \N__3652\,
            I => \N__3642\
        );

    \I__471\ : InMux
    port map (
            O => \N__3651\,
            I => \N__3642\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3642\,
            I => \N__3636\
        );

    \I__469\ : InMux
    port map (
            O => \N__3641\,
            I => \N__3629\
        );

    \I__468\ : InMux
    port map (
            O => \N__3640\,
            I => \N__3629\
        );

    \I__467\ : InMux
    port map (
            O => \N__3639\,
            I => \N__3629\
        );

    \I__466\ : Odrv4
    port map (
            O => \N__3636\,
            I => \fsm_ctrl_inst1.counter_stat12_i_0\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3629\,
            I => \fsm_ctrl_inst1.counter_stat12_i_0\
        );

    \I__464\ : InMux
    port map (
            O => \N__3624\,
            I => \N__3621\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__3621\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_0\
        );

    \I__462\ : InMux
    port map (
            O => \N__3618\,
            I => \N__3615\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__3615\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_1\
        );

    \I__460\ : InMux
    port map (
            O => \N__3612\,
            I => \N__3609\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3609\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_2\
        );

    \I__458\ : InMux
    port map (
            O => \N__3606\,
            I => \N__3603\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3603\,
            I => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_3\
        );

    \I__456\ : InMux
    port map (
            O => \N__3600\,
            I => \N__3597\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__3597\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_56\
        );

    \I__454\ : InMux
    port map (
            O => \N__3594\,
            I => \N__3591\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3591\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_57\
        );

    \I__452\ : InMux
    port map (
            O => \N__3588\,
            I => \N__3585\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__3585\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_54\
        );

    \I__450\ : InMux
    port map (
            O => \N__3582\,
            I => \N__3579\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__3579\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_55\
        );

    \I__448\ : InMux
    port map (
            O => \N__3576\,
            I => \N__3573\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__3573\,
            I => \N__3570\
        );

    \I__446\ : Odrv12
    port map (
            O => \N__3570\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_23\
        );

    \I__445\ : InMux
    port map (
            O => \N__3567\,
            I => \N__3564\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__3564\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_24\
        );

    \I__443\ : InMux
    port map (
            O => \N__3561\,
            I => \N__3558\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__3558\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_48\
        );

    \I__441\ : InMux
    port map (
            O => \N__3555\,
            I => \N__3552\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__3552\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_49\
        );

    \I__439\ : InMux
    port map (
            O => \N__3549\,
            I => \N__3546\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__3546\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_45\
        );

    \I__437\ : InMux
    port map (
            O => \N__3543\,
            I => \N__3540\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3540\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_43\
        );

    \I__435\ : CascadeMux
    port map (
            O => \N__3537\,
            I => \fsm_ctrl_inst1.current_state_ns_i_i_a2_0_5_1_cascade_\
        );

    \I__434\ : IoInMux
    port map (
            O => \N__3534\,
            I => \N__3531\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__3531\,
            I => \N__3528\
        );

    \I__432\ : Span4Mux_s2_h
    port map (
            O => \N__3528\,
            I => \N__3525\
        );

    \I__431\ : Odrv4
    port map (
            O => \N__3525\,
            I => \fsm_ctrl_inst1.current_state_i_0\
        );

    \I__430\ : InMux
    port map (
            O => \N__3522\,
            I => \N__3518\
        );

    \I__429\ : InMux
    port map (
            O => \N__3521\,
            I => \N__3515\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3518\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_0\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3515\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_0\
        );

    \I__426\ : InMux
    port map (
            O => \N__3510\,
            I => \bfn_3_20_0_\
        );

    \I__425\ : InMux
    port map (
            O => \N__3507\,
            I => \N__3500\
        );

    \I__424\ : InMux
    port map (
            O => \N__3506\,
            I => \N__3500\
        );

    \I__423\ : InMux
    port map (
            O => \N__3505\,
            I => \N__3497\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__3500\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_1\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3497\,
            I => \fsm_ctrl_inst1.counter_idleZ0Z_1\
        );

    \I__420\ : InMux
    port map (
            O => \N__3492\,
            I => \fsm_ctrl_inst1.counter_idle_cry_0\
        );

    \I__419\ : InMux
    port map (
            O => \N__3489\,
            I => \fsm_ctrl_inst1.counter_idle_cry_1\
        );

    \I__418\ : InMux
    port map (
            O => \N__3486\,
            I => \fsm_ctrl_inst1.counter_idle_cry_2\
        );

    \I__417\ : InMux
    port map (
            O => \N__3483\,
            I => \fsm_ctrl_inst1.counter_idle_cry_3\
        );

    \I__416\ : CEMux
    port map (
            O => \N__3480\,
            I => \N__3477\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__3477\,
            I => \N__3474\
        );

    \I__414\ : Odrv4
    port map (
            O => \N__3474\,
            I => \fsm_ctrl_inst1.counter_idlee_0_i\
        );

    \I__413\ : InMux
    port map (
            O => \N__3471\,
            I => \fsm_ctrl_inst1.counter_stat_cry_1\
        );

    \I__412\ : InMux
    port map (
            O => \N__3468\,
            I => \fsm_ctrl_inst1.counter_stat_cry_2\
        );

    \I__411\ : InMux
    port map (
            O => \N__3465\,
            I => \fsm_ctrl_inst1.counter_stat_cry_3\
        );

    \I__410\ : InMux
    port map (
            O => \N__3462\,
            I => \fsm_ctrl_inst1.counter_stat_cry_4\
        );

    \I__409\ : InMux
    port map (
            O => \N__3459\,
            I => \fsm_ctrl_inst1.counter_stat_cry_5\
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__3456\,
            I => \fsm_ctrl_inst1.current_state_ns_0_i_0_1_0_cascade_\
        );

    \I__407\ : CascadeMux
    port map (
            O => \N__3453\,
            I => \N__3449\
        );

    \I__406\ : InMux
    port map (
            O => \N__3452\,
            I => \N__3446\
        );

    \I__405\ : InMux
    port map (
            O => \N__3449\,
            I => \N__3443\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__3446\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_1\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__3443\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_1\
        );

    \I__402\ : InMux
    port map (
            O => \N__3438\,
            I => \N__3434\
        );

    \I__401\ : InMux
    port map (
            O => \N__3437\,
            I => \N__3431\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__3434\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_0\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__3431\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_0\
        );

    \I__398\ : InMux
    port map (
            O => \N__3426\,
            I => \N__3422\
        );

    \I__397\ : InMux
    port map (
            O => \N__3425\,
            I => \N__3419\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__3422\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_2\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__3419\,
            I => \fsm_ctrl_inst1.counter_statZ0Z_2\
        );

    \I__394\ : CascadeMux
    port map (
            O => \N__3414\,
            I => \fsm_ctrl_inst1.current_state_ns_i_i_a2_0_4_1_cascade_\
        );

    \I__393\ : InMux
    port map (
            O => \N__3411\,
            I => \N__3408\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__3408\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_16\
        );

    \I__391\ : InMux
    port map (
            O => \N__3405\,
            I => \N__3402\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3402\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_42\
        );

    \I__389\ : InMux
    port map (
            O => \N__3399\,
            I => \N__3396\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__3396\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_19\
        );

    \I__387\ : InMux
    port map (
            O => \N__3393\,
            I => \N__3390\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__3390\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_17\
        );

    \I__385\ : InMux
    port map (
            O => \N__3387\,
            I => \N__3384\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__3384\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_18\
        );

    \I__383\ : InMux
    port map (
            O => \N__3381\,
            I => \N__3378\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3378\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_20\
        );

    \I__381\ : InMux
    port map (
            O => \N__3375\,
            I => \N__3372\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__3372\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_21\
        );

    \I__379\ : InMux
    port map (
            O => \N__3369\,
            I => \N__3366\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__3366\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_22\
        );

    \I__377\ : InMux
    port map (
            O => \N__3363\,
            I => \bfn_3_18_0_\
        );

    \I__376\ : InMux
    port map (
            O => \N__3360\,
            I => \fsm_ctrl_inst1.counter_stat_cry_0\
        );

    \I__375\ : InMux
    port map (
            O => \N__3357\,
            I => \N__3354\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__3354\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_29\
        );

    \I__373\ : InMux
    port map (
            O => \N__3351\,
            I => \N__3348\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__3348\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_25\
        );

    \I__371\ : InMux
    port map (
            O => \N__3345\,
            I => \N__3342\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__3342\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_26\
        );

    \I__369\ : InMux
    port map (
            O => \N__3339\,
            I => \N__3336\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__3336\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_5\
        );

    \I__367\ : InMux
    port map (
            O => \N__3333\,
            I => \N__3330\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__3330\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_6\
        );

    \I__365\ : InMux
    port map (
            O => \N__3327\,
            I => \N__3324\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__3324\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_7\
        );

    \I__363\ : InMux
    port map (
            O => \N__3321\,
            I => \N__3318\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__3318\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_27\
        );

    \I__361\ : InMux
    port map (
            O => \N__3315\,
            I => \N__3312\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__3312\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_28\
        );

    \I__359\ : InMux
    port map (
            O => \N__3309\,
            I => \N__3306\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3306\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_58\
        );

    \I__357\ : InMux
    port map (
            O => \N__3303\,
            I => \N__3300\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__3300\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_32\
        );

    \I__355\ : InMux
    port map (
            O => \N__3297\,
            I => \N__3294\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__3294\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_10\
        );

    \I__353\ : InMux
    port map (
            O => \N__3291\,
            I => \N__3288\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__3288\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_9\
        );

    \I__351\ : InMux
    port map (
            O => \N__3285\,
            I => \N__3282\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__3282\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_31\
        );

    \I__349\ : InMux
    port map (
            O => \N__3279\,
            I => \N__3276\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__3276\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_3\
        );

    \I__347\ : InMux
    port map (
            O => \N__3273\,
            I => \N__3270\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__3270\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_4\
        );

    \I__345\ : InMux
    port map (
            O => \N__3267\,
            I => \N__3264\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__3264\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_59\
        );

    \I__343\ : InMux
    port map (
            O => \N__3261\,
            I => \N__3258\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__3258\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_30\
        );

    \I__341\ : InMux
    port map (
            O => \N__3255\,
            I => \N__3252\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__3252\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_8\
        );

    \I__339\ : InMux
    port map (
            O => \N__3249\,
            I => \N__3246\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__3246\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_36\
        );

    \I__337\ : InMux
    port map (
            O => \N__3243\,
            I => \N__3240\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__3240\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_37\
        );

    \I__335\ : InMux
    port map (
            O => \N__3237\,
            I => \N__3234\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__3234\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_38\
        );

    \I__333\ : InMux
    port map (
            O => \N__3231\,
            I => \N__3228\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__3228\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_1\
        );

    \I__331\ : InMux
    port map (
            O => \N__3225\,
            I => \N__3222\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__3222\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_0\
        );

    \I__329\ : InMux
    port map (
            O => \N__3219\,
            I => \N__3216\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__3216\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_11\
        );

    \I__327\ : InMux
    port map (
            O => \N__3213\,
            I => \N__3210\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__3210\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_62\
        );

    \I__325\ : InMux
    port map (
            O => \N__3207\,
            I => \N__3204\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__3204\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_60\
        );

    \I__323\ : InMux
    port map (
            O => \N__3201\,
            I => \N__3198\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__3198\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_61\
        );

    \I__321\ : InMux
    port map (
            O => \N__3195\,
            I => \N__3192\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__3192\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_82\
        );

    \I__319\ : InMux
    port map (
            O => \N__3189\,
            I => \N__3186\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__3186\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_67\
        );

    \I__317\ : InMux
    port map (
            O => \N__3183\,
            I => \N__3180\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__3180\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_14\
        );

    \I__315\ : InMux
    port map (
            O => \N__3177\,
            I => \N__3174\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__3174\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_15\
        );

    \I__313\ : InMux
    port map (
            O => \N__3171\,
            I => \N__3168\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__3168\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_13\
        );

    \I__311\ : InMux
    port map (
            O => \N__3165\,
            I => \N__3162\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__3162\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_63\
        );

    \I__309\ : InMux
    port map (
            O => \N__3159\,
            I => \N__3156\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__3156\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_40\
        );

    \I__307\ : InMux
    port map (
            O => \N__3153\,
            I => \N__3150\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__3150\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_41\
        );

    \I__305\ : InMux
    port map (
            O => \N__3147\,
            I => \N__3144\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__3144\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_12\
        );

    \I__303\ : InMux
    port map (
            O => \N__3141\,
            I => \N__3138\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__3138\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_39\
        );

    \I__301\ : InMux
    port map (
            O => \N__3135\,
            I => \N__3132\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__3132\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_33\
        );

    \I__299\ : InMux
    port map (
            O => \N__3129\,
            I => \N__3126\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__3126\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_80\
        );

    \I__297\ : InMux
    port map (
            O => \N__3123\,
            I => \N__3120\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__3120\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_81\
        );

    \I__295\ : InMux
    port map (
            O => \N__3117\,
            I => \N__3114\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__3114\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_2\
        );

    \I__293\ : InMux
    port map (
            O => \N__3111\,
            I => \N__3108\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__3108\,
            I => \N__3105\
        );

    \I__291\ : Odrv4
    port map (
            O => \N__3105\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_70\
        );

    \I__290\ : InMux
    port map (
            O => \N__3102\,
            I => \N__3099\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__3099\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_68\
        );

    \I__288\ : InMux
    port map (
            O => \N__3096\,
            I => \N__3093\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__3093\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_69\
        );

    \I__286\ : InMux
    port map (
            O => \N__3090\,
            I => \N__3087\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__3087\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_66\
        );

    \I__284\ : InMux
    port map (
            O => \N__3084\,
            I => \N__3081\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__3081\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_73\
        );

    \I__282\ : InMux
    port map (
            O => \N__3078\,
            I => \N__3075\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__3075\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_74\
        );

    \I__280\ : InMux
    port map (
            O => \N__3072\,
            I => \N__3069\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__3069\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_75\
        );

    \I__278\ : InMux
    port map (
            O => \N__3066\,
            I => \N__3063\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__3063\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_35\
        );

    \I__276\ : InMux
    port map (
            O => \N__3060\,
            I => \N__3057\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__3057\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_79\
        );

    \I__274\ : InMux
    port map (
            O => \N__3054\,
            I => \N__3051\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__3051\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_78\
        );

    \I__272\ : InMux
    port map (
            O => \N__3048\,
            I => \N__3045\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__3045\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_76\
        );

    \I__270\ : InMux
    port map (
            O => \N__3042\,
            I => \N__3039\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__3039\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_77\
        );

    \I__268\ : InMux
    port map (
            O => \N__3036\,
            I => \N__3033\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__3033\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_34\
        );

    \I__266\ : InMux
    port map (
            O => \N__3030\,
            I => \N__3027\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__3027\,
            I => \RST_N_c\
        );

    \I__264\ : IoInMux
    port map (
            O => \N__3024\,
            I => \N__3021\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__3021\,
            I => \RST_N_c_i\
        );

    \I__262\ : InMux
    port map (
            O => \N__3018\,
            I => \N__3015\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__3015\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_72\
        );

    \I__260\ : InMux
    port map (
            O => \N__3012\,
            I => \N__3009\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__3009\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_71\
        );

    \I__258\ : InMux
    port map (
            O => \N__3006\,
            I => \N__3003\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__3003\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_64\
        );

    \I__256\ : InMux
    port map (
            O => \N__3000\,
            I => \N__2997\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2997\,
            I => \fsm_ctrl_inst1.bit_sequence_statZ0Z_65\
        );

    \IN_MUX_bfv_3_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_18_0_\
        );

    \IN_MUX_bfv_3_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_20_0_\
        );

    \fsm_ctrl_inst1.SEL_RNIQ5L_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4638\,
            GLOBALBUFFEROUTPUT => \SEL_REG_i_g\
        );

    \fsm_ctrl_inst1.current_state_RNI1GR8_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3534\,
            GLOBALBUFFEROUTPUT => \fsm_ctrl_inst1.current_state_i_g_0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \RST_N_ibuf_RNIBJGC_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3024\,
            GLOBALBUFFEROUTPUT => \RST_N_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \RST_N_ibuf_RNIBJGC_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3030\,
            lcout => \RST_N_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_72_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3012\,
            in2 => \_gnd_net_\,
            in3 => \N__4333\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5710\,
            ce => \N__4388\,
            sr => \N__5434\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_65_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4330\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3006\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5710\,
            ce => \N__4388\,
            sr => \N__5434\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_73_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3018\,
            in2 => \_gnd_net_\,
            in3 => \N__4334\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5710\,
            ce => \N__4388\,
            sr => \N__5434\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_71_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4332\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3111\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5710\,
            ce => \N__4388\,
            sr => \N__5434\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_64_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3165\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4329\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5710\,
            ce => \N__4388\,
            sr => \N__5434\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_66_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4331\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3000\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5710\,
            ce => \N__4388\,
            sr => \N__5434\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_76_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3072\,
            in2 => \_gnd_net_\,
            in3 => \N__4326\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5712\,
            ce => \N__4390\,
            sr => \N__5435\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_74_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__3084\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4324\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5712\,
            ce => \N__4390\,
            sr => \N__5435\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_75_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4325\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3078\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5712\,
            ce => \N__4390\,
            sr => \N__5435\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_36_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3066\,
            in2 => \_gnd_net_\,
            in3 => \N__4323\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5712\,
            ce => \N__4390\,
            sr => \N__5435\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_35_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3036\,
            in2 => \_gnd_net_\,
            in3 => \N__4322\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5712\,
            ce => \N__4390\,
            sr => \N__5435\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_80_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4287\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3060\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5714\,
            ce => \N__4392\,
            sr => \N__5437\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_79_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4286\,
            in2 => \_gnd_net_\,
            in3 => \N__3054\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5714\,
            ce => \N__4392\,
            sr => \N__5437\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_78_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4285\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3042\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5714\,
            ce => \N__4392\,
            sr => \N__5437\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_77_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1011101110111011"
        )
    port map (
            in0 => \N__3048\,
            in1 => \N__4284\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5714\,
            ce => \N__4392\,
            sr => \N__5437\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_34_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4283\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3135\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5714\,
            ce => \N__4392\,
            sr => \N__5437\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_33_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4282\,
            in2 => \_gnd_net_\,
            in3 => \N__3303\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5714\,
            ce => \N__4392\,
            sr => \N__5437\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_81_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4288\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3129\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5714\,
            ce => \N__4392\,
            sr => \N__5437\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_82_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4289\,
            in2 => \_gnd_net_\,
            in3 => \N__3123\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5714\,
            ce => \N__4392\,
            sr => \N__5437\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_3_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4328\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3117\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5717\,
            ce => \N__4395\,
            sr => \N__5440\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_2_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3231\,
            in2 => \_gnd_net_\,
            in3 => \N__4327\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5717\,
            ce => \N__4395\,
            sr => \N__5440\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_70_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4254\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3096\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5711\,
            ce => \N__4389\,
            sr => \N__5436\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_68_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3189\,
            in2 => \_gnd_net_\,
            in3 => \N__4252\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5711\,
            ce => \N__4389\,
            sr => \N__5436\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_69_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4253\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3102\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5711\,
            ce => \N__4389\,
            sr => \N__5436\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_14_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3171\,
            in2 => \_gnd_net_\,
            in3 => \N__4248\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5711\,
            ce => \N__4389\,
            sr => \N__5436\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_67_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4251\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3090\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5711\,
            ce => \N__4389\,
            sr => \N__5436\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_16_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3177\,
            in2 => \_gnd_net_\,
            in3 => \N__4250\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5711\,
            ce => \N__4389\,
            sr => \N__5436\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_15_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4249\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3183\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5711\,
            ce => \N__4389\,
            sr => \N__5436\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_13_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3147\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4247\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5711\,
            ce => \N__4389\,
            sr => \N__5436\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_63_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3213\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4221\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5715\,
            ce => \N__4393\,
            sr => \N__5438\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_40_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4218\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3141\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5715\,
            ce => \N__4393\,
            sr => \N__5438\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_41_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3159\,
            in2 => \_gnd_net_\,
            in3 => \N__4219\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5715\,
            ce => \N__4393\,
            sr => \N__5438\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_42_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4220\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3153\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5715\,
            ce => \N__4393\,
            sr => \N__5438\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_12_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3219\,
            in2 => \_gnd_net_\,
            in3 => \N__4214\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5715\,
            ce => \N__4393\,
            sr => \N__5438\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_39_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4217\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3237\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5715\,
            ce => \N__4393\,
            sr => \N__5438\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_37_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3249\,
            in2 => \_gnd_net_\,
            in3 => \N__4215\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5715\,
            ce => \N__4393\,
            sr => \N__5438\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_38_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4216\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3243\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5715\,
            ce => \N__4393\,
            sr => \N__5438\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_1_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3225\,
            in2 => \_gnd_net_\,
            in3 => \N__4094\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5718\,
            ce => \N__4396\,
            sr => \N__5441\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_60_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4096\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3267\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5718\,
            ce => \N__4396\,
            sr => \N__5441\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_0_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4092\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5718\,
            ce => \N__4396\,
            sr => \N__5441\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_11_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__4093\,
            in1 => \N__3297\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5718\,
            ce => \N__4396\,
            sr => \N__5441\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_62_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3201\,
            in2 => \_gnd_net_\,
            in3 => \N__4098\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5718\,
            ce => \N__4396\,
            sr => \N__5441\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_61_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4097\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3207\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5718\,
            ce => \N__4396\,
            sr => \N__5441\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_83_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3195\,
            in2 => \_gnd_net_\,
            in3 => \N__4099\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5718\,
            ce => \N__4396\,
            sr => \N__5441\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_32_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4095\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3285\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5718\,
            ce => \N__4396\,
            sr => \N__5441\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_10_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3291\,
            in2 => \_gnd_net_\,
            in3 => \N__4206\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5720\,
            ce => \N__4397\,
            sr => \N__5444\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_9_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4213\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3255\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5720\,
            ce => \N__4397\,
            sr => \N__5444\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_31_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3261\,
            in2 => \_gnd_net_\,
            in3 => \N__4208\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5720\,
            ce => \N__4397\,
            sr => \N__5444\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_5_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4211\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3273\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5720\,
            ce => \N__4397\,
            sr => \N__5444\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_4_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3279\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4209\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5720\,
            ce => \N__4397\,
            sr => \N__5444\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_59_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4210\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3309\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5720\,
            ce => \N__4397\,
            sr => \N__5444\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_30_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3357\,
            in2 => \_gnd_net_\,
            in3 => \N__4207\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5720\,
            ce => \N__4397\,
            sr => \N__5444\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_8_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4212\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3327\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5720\,
            ce => \N__4397\,
            sr => \N__5444\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_26_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3351\,
            in2 => \_gnd_net_\,
            in3 => \N__4264\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5723\,
            ce => \N__4398\,
            sr => \N__5447\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_29_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4267\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3315\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5723\,
            ce => \N__4398\,
            sr => \N__5447\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_25_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3567\,
            in2 => \_gnd_net_\,
            in3 => \N__4263\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5723\,
            ce => \N__4398\,
            sr => \N__5447\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_27_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4265\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3345\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5723\,
            ce => \N__4398\,
            sr => \N__5447\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_6_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3339\,
            in2 => \_gnd_net_\,
            in3 => \N__4269\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5723\,
            ce => \N__4398\,
            sr => \N__5447\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_7_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4270\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3333\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5723\,
            ce => \N__4398\,
            sr => \N__5447\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_28_LC_2_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3321\,
            in2 => \_gnd_net_\,
            in3 => \N__4266\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5723\,
            ce => \N__4398\,
            sr => \N__5447\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_58_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4268\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3594\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5723\,
            ce => \N__4398\,
            sr => \N__5447\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_19_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4241\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3387\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5713\,
            ce => \N__4391\,
            sr => \N__5439\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_17_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3411\,
            in2 => \_gnd_net_\,
            in3 => \N__4239\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5713\,
            ce => \N__4391\,
            sr => \N__5439\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_23_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4245\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3369\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5713\,
            ce => \N__4391\,
            sr => \N__5439\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_43_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3405\,
            in2 => \_gnd_net_\,
            in3 => \N__4246\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5713\,
            ce => \N__4391\,
            sr => \N__5439\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_20_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4242\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3399\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5713\,
            ce => \N__4391\,
            sr => \N__5439\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_18_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3393\,
            in2 => \_gnd_net_\,
            in3 => \N__4240\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5713\,
            ce => \N__4391\,
            sr => \N__5439\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_21_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4243\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3381\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5713\,
            ce => \N__4391\,
            sr => \N__5439\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_22_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3375\,
            in2 => \_gnd_net_\,
            in3 => \N__4244\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5713\,
            ce => \N__4391\,
            sr => \N__5439\
        );

    \fsm_ctrl_inst1.counter_stat_0_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3651\,
            in1 => \N__3438\,
            in2 => \_gnd_net_\,
            in3 => \N__3363\,
            lcout => \fsm_ctrl_inst1.counter_statZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_3_18_0_\,
            carryout => \fsm_ctrl_inst1.counter_stat_cry_0\,
            clk => \N__5719\,
            ce => \N__3834\,
            sr => \N__5442\
        );

    \fsm_ctrl_inst1.counter_stat_1_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3639\,
            in1 => \N__3452\,
            in2 => \_gnd_net_\,
            in3 => \N__3360\,
            lcout => \fsm_ctrl_inst1.counter_statZ0Z_1\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_stat_cry_0\,
            carryout => \fsm_ctrl_inst1.counter_stat_cry_1\,
            clk => \N__5719\,
            ce => \N__3834\,
            sr => \N__5442\
        );

    \fsm_ctrl_inst1.counter_stat_2_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3652\,
            in1 => \N__3425\,
            in2 => \_gnd_net_\,
            in3 => \N__3471\,
            lcout => \fsm_ctrl_inst1.counter_statZ0Z_2\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_stat_cry_1\,
            carryout => \fsm_ctrl_inst1.counter_stat_cry_2\,
            clk => \N__5719\,
            ce => \N__3834\,
            sr => \N__5442\
        );

    \fsm_ctrl_inst1.counter_stat_3_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3640\,
            in1 => \N__3716\,
            in2 => \_gnd_net_\,
            in3 => \N__3468\,
            lcout => \fsm_ctrl_inst1.counter_statZ0Z_3\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_stat_cry_2\,
            carryout => \fsm_ctrl_inst1.counter_stat_cry_3\,
            clk => \N__5719\,
            ce => \N__3834\,
            sr => \N__5442\
        );

    \fsm_ctrl_inst1.counter_stat_4_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3653\,
            in1 => \N__3736\,
            in2 => \_gnd_net_\,
            in3 => \N__3465\,
            lcout => \fsm_ctrl_inst1.counter_statZ0Z_4\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_stat_cry_3\,
            carryout => \fsm_ctrl_inst1.counter_stat_cry_4\,
            clk => \N__5719\,
            ce => \N__3834\,
            sr => \N__5442\
        );

    \fsm_ctrl_inst1.counter_stat_5_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3641\,
            in1 => \N__3695\,
            in2 => \_gnd_net_\,
            in3 => \N__3462\,
            lcout => \fsm_ctrl_inst1.counter_statZ0Z_5\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_stat_cry_4\,
            carryout => \fsm_ctrl_inst1.counter_stat_cry_5\,
            clk => \N__5719\,
            ce => \N__3834\,
            sr => \N__5442\
        );

    \fsm_ctrl_inst1.counter_stat_6_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3654\,
            in1 => \N__3675\,
            in2 => \_gnd_net_\,
            in3 => \N__3459\,
            lcout => \fsm_ctrl_inst1.counter_statZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5719\,
            ce => \N__3834\,
            sr => \N__5442\
        );

    \fsm_ctrl_inst1.current_state_RNO_0_0_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__3522\,
            in1 => \N__3506\,
            in2 => \_gnd_net_\,
            in3 => \N__4087\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.current_state_ns_0_i_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.current_state_0_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__4702\,
            in1 => \N__4505\,
            in2 => \N__3456\,
            in3 => \N__3765\,
            lcout => \fsm_ctrl_inst1.current_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5721\,
            ce => 'H',
            sr => \N__5445\
        );

    \fsm_ctrl_inst1.current_state_RNO_1_1_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__3674\,
            in1 => \N__3694\,
            in2 => \N__3453\,
            in3 => \N__3437\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.current_state_ns_i_i_a2_0_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.current_state_RNO_0_1_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__3426\,
            in1 => \N__3737\,
            in2 => \N__3414\,
            in3 => \N__3717\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.current_state_ns_i_i_a2_0_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.current_state_1_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001110100001100"
        )
    port map (
            in0 => \N__4506\,
            in1 => \N__4091\,
            in2 => \N__3537\,
            in3 => \N__4703\,
            lcout => \fsm_ctrl_inst1.current_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5721\,
            ce => 'H',
            sr => \N__5445\
        );

    \fsm_ctrl_inst1.current_state_RNI1GR8_0_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4701\,
            lcout => \fsm_ctrl_inst1.current_state_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_RNIPMA12_1_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__3507\,
            in1 => \N__4710\,
            in2 => \N__4238\,
            in3 => \N__3764\,
            lcout => \fsm_ctrl_inst1.counter_idlee_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_0_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3829\,
            in1 => \N__3521\,
            in2 => \_gnd_net_\,
            in3 => \N__3510\,
            lcout => \fsm_ctrl_inst1.counter_idleZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_3_20_0_\,
            carryout => \fsm_ctrl_inst1.counter_idle_cry_0\,
            clk => \N__5724\,
            ce => \N__3480\,
            sr => \N__5448\
        );

    \fsm_ctrl_inst1.counter_idle_1_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3826\,
            in1 => \N__3505\,
            in2 => \_gnd_net_\,
            in3 => \N__3492\,
            lcout => \fsm_ctrl_inst1.counter_idleZ0Z_1\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_idle_cry_0\,
            carryout => \fsm_ctrl_inst1.counter_idle_cry_1\,
            clk => \N__5724\,
            ce => \N__3480\,
            sr => \N__5448\
        );

    \fsm_ctrl_inst1.counter_idle_2_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3830\,
            in1 => \N__3789\,
            in2 => \_gnd_net_\,
            in3 => \N__3489\,
            lcout => \fsm_ctrl_inst1.counter_idleZ0Z_2\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_idle_cry_1\,
            carryout => \fsm_ctrl_inst1.counter_idle_cry_2\,
            clk => \N__5724\,
            ce => \N__3480\,
            sr => \N__5448\
        );

    \fsm_ctrl_inst1.counter_idle_3_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3827\,
            in1 => \N__3801\,
            in2 => \_gnd_net_\,
            in3 => \N__3486\,
            lcout => \fsm_ctrl_inst1.counter_idleZ0Z_3\,
            ltout => OPEN,
            carryin => \fsm_ctrl_inst1.counter_idle_cry_2\,
            carryout => \fsm_ctrl_inst1.counter_idle_cry_3\,
            clk => \N__5724\,
            ce => \N__3480\,
            sr => \N__5448\
        );

    \fsm_ctrl_inst1.counter_idle_4_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__3777\,
            in1 => \N__3828\,
            in2 => \_gnd_net_\,
            in3 => \N__3483\,
            lcout => \fsm_ctrl_inst1.counter_idleZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5724\,
            ce => \N__3480\,
            sr => \N__5448\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_50_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3555\,
            in2 => \_gnd_net_\,
            in3 => \N__4258\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5726\,
            ce => \N__4399\,
            sr => \N__5450\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_56_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4261\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3582\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5726\,
            ce => \N__4399\,
            sr => \N__5450\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_57_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3600\,
            in2 => \_gnd_net_\,
            in3 => \N__4262\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5726\,
            ce => \N__4399\,
            sr => \N__5450\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_48_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4256\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3894\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5726\,
            ce => \N__4399\,
            sr => \N__5450\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_54_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3888\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4259\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5726\,
            ce => \N__4399\,
            sr => \N__5450\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_55_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4260\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3588\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5726\,
            ce => \N__4399\,
            sr => \N__5450\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_24_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3576\,
            in2 => \_gnd_net_\,
            in3 => \N__4255\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5726\,
            ce => \N__4399\,
            sr => \N__5450\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_49_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4257\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3561\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5726\,
            ce => \N__4399\,
            sr => \N__5450\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_46_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3549\,
            in2 => \_gnd_net_\,
            in3 => \N__4317\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5716\,
            ce => \N__4394\,
            sr => \N__5443\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_45_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4316\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3744\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5716\,
            ce => \N__4394\,
            sr => \N__5443\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_44_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3543\,
            in2 => \_gnd_net_\,
            in3 => \N__4315\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5716\,
            ce => \N__4394\,
            sr => \N__5443\
        );

    \fsm_ctrl_inst1.counter_stat_RNIML9_6_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__3738\,
            in1 => \N__3715\,
            in2 => \N__3699\,
            in3 => \N__3673\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.counter_stat_RNIML9Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.current_state_RNIO659_1_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__3864\,
            in1 => \_gnd_net_\,
            in2 => \N__3657\,
            in3 => \N__4084\,
            lcout => \fsm_ctrl_inst1.counter_stat12_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.current_state_RNI2HR8_1_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4085\,
            lcout => \fsm_ctrl_inst1.current_state_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.bit_sequence_din_0_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4727\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5722\,
            ce => \N__3919\,
            sr => \N__5446\
        );

    \fsm_ctrl_inst1.bit_sequence_din_1_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4725\,
            in2 => \_gnd_net_\,
            in3 => \N__3624\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5722\,
            ce => \N__3919\,
            sr => \N__5446\
        );

    \fsm_ctrl_inst1.bit_sequence_din_2_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__4728\,
            in1 => \N__3618\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5722\,
            ce => \N__3919\,
            sr => \N__5446\
        );

    \fsm_ctrl_inst1.bit_sequence_din_3_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4726\,
            in2 => \_gnd_net_\,
            in3 => \N__3612\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5722\,
            ce => \N__3919\,
            sr => \N__5446\
        );

    \fsm_ctrl_inst1.bit_sequence_din_4_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4705\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3606\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5725\,
            ce => \N__3920\,
            sr => \N__5449\
        );

    \fsm_ctrl_inst1.bit_sequence_din_5_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3858\,
            in2 => \_gnd_net_\,
            in3 => \N__4708\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5725\,
            ce => \N__3920\,
            sr => \N__5449\
        );

    \fsm_ctrl_inst1.bit_sequence_din_6_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4706\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3852\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5725\,
            ce => \N__3920\,
            sr => \N__5449\
        );

    \fsm_ctrl_inst1.bit_sequence_din_7_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3846\,
            in2 => \_gnd_net_\,
            in3 => \N__4709\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5725\,
            ce => \N__3920\,
            sr => \N__5449\
        );

    \fsm_ctrl_inst1.bit_sequence_din_8_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4707\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3840\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5725\,
            ce => \N__3920\,
            sr => \N__5449\
        );

    \fsm_ctrl_inst1.current_state_RNI31NH_0_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4086\,
            in2 => \_gnd_net_\,
            in3 => \N__4704\,
            lcout => \fsm_ctrl_inst1.counter_state_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_idle_RNIQPM31_4_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3800\,
            in1 => \N__3788\,
            in2 => \_gnd_net_\,
            in3 => \N__3776\,
            lcout => \fsm_ctrl_inst1.N_127_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.bit_sequence_din_10_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3930\,
            in2 => \_gnd_net_\,
            in3 => \N__4721\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5727\,
            ce => \N__3924\,
            sr => \N__5451\
        );

    \fsm_ctrl_inst1.bit_sequence_din_11_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4718\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3756\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5727\,
            ce => \N__3924\,
            sr => \N__5451\
        );

    \fsm_ctrl_inst1.bit_sequence_din_12_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3750\,
            in2 => \_gnd_net_\,
            in3 => \N__4722\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5727\,
            ce => \N__3924\,
            sr => \N__5451\
        );

    \fsm_ctrl_inst1.bit_sequence_din_13_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4719\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3957\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5727\,
            ce => \N__3924\,
            sr => \N__5451\
        );

    \fsm_ctrl_inst1.bit_sequence_din_14_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3951\,
            in2 => \_gnd_net_\,
            in3 => \N__4723\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5727\,
            ce => \N__3924\,
            sr => \N__5451\
        );

    \fsm_ctrl_inst1.bit_sequence_din_15_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4720\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3945\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5727\,
            ce => \N__3924\,
            sr => \N__5451\
        );

    \fsm_ctrl_inst1.bit_sequence_din_9_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3939\,
            in2 => \_gnd_net_\,
            in3 => \N__4724\,
            lcout => \fsm_ctrl_inst1.bit_sequence_dinZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5727\,
            ce => \N__3924\,
            sr => \N__5451\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_47_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3903\,
            in2 => \_gnd_net_\,
            in3 => \N__4318\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5729\,
            ce => \N__4401\,
            sr => \N__5453\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_53_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4321\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3882\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5729\,
            ce => \N__4401\,
            sr => \N__5453\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_52_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3870\,
            in2 => \_gnd_net_\,
            in3 => \N__4320\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5729\,
            ce => \N__4401\,
            sr => \N__5453\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_51_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3876\,
            in2 => \_gnd_net_\,
            in3 => \N__4319\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5729\,
            ce => \N__4401\,
            sr => \N__5453\
        );

    \CONSTANT_ONE_LUT4_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_85_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4419\,
            in2 => \_gnd_net_\,
            in3 => \N__4312\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5728\,
            ce => \N__4400\,
            sr => \N__5452\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_87_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4407\,
            in2 => \_gnd_net_\,
            in3 => \N__4314\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5728\,
            ce => \N__4400\,
            sr => \N__5452\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_84_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4428\,
            in2 => \_gnd_net_\,
            in3 => \N__4311\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5728\,
            ce => \N__4400\,
            sr => \N__5452\
        );

    \fsm_ctrl_inst1.bit_sequence_stat_86_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4413\,
            in2 => \_gnd_net_\,
            in3 => \N__4313\,
            lcout => \fsm_ctrl_inst1.bit_sequence_statZ0Z_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5728\,
            ce => \N__4400\,
            sr => \N__5452\
        );

    \fsm_ctrl_inst1.MOSI_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__4744\,
            in1 => \N__4353\,
            in2 => \N__4347\,
            in3 => \N__4335\,
            lcout => \MOSI\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5730\,
            ce => 'H',
            sr => \N__5454\
        );

    \fsm_ctrl_inst1.counter_din_0_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4466\,
            in2 => \_gnd_net_\,
            in3 => \N__4745\,
            lcout => \fsm_ctrl_inst1.counter_dinZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5730\,
            ce => 'H',
            sr => \N__5454\
        );

    \config_register_latched_dec_inst1.DYNSR_1_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4575\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5731\,
            ce => \N__4810\,
            sr => \N__5455\
        );

    \config_register_latched_dec_inst1.DYNSR_4_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4563\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5731\,
            ce => \N__4810\,
            sr => \N__5455\
        );

    \config_register_latched_dec_inst1.DYNSR_2_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3963\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5731\,
            ce => \N__4810\,
            sr => \N__5455\
        );

    \config_register_latched_dec_inst1.DYNSR_0_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4553\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5731\,
            ce => \N__4810\,
            sr => \N__5455\
        );

    \config_register_latched_dec_inst1.DYNSR_3_LC_5_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4569\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5731\,
            ce => \N__4810\,
            sr => \N__5455\
        );

    \config_register_latched_dec_inst1.STATSR_0_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4557\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5734\,
            ce => \N__5589\,
            sr => \N__5458\
        );

    \config_register_latched_dec_inst1.DYNSR_RNIQ2U9_15_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__4805\,
            in1 => \N__4977\,
            in2 => \_gnd_net_\,
            in3 => \N__4863\,
            lcout => \SDO_signal_out_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_din_RNO_0_3_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__4441\,
            in1 => \N__4517\,
            in2 => \N__4484\,
            in3 => \N__4461\,
            lcout => OPEN,
            ltout => \fsm_ctrl_inst1.counter_din_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_din_3_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4747\,
            in2 => \N__4521\,
            in3 => \N__4496\,
            lcout => \fsm_ctrl_inst1.counter_dinZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5732\,
            ce => 'H',
            sr => \N__5456\
        );

    \fsm_ctrl_inst1.counter_din_RNI6L3H1_3_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__4460\,
            in1 => \N__4477\,
            in2 => \N__4518\,
            in3 => \N__4440\,
            lcout => \fsm_ctrl_inst1.counter_din_RNI6L3H1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fsm_ctrl_inst1.counter_din_2_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100000000000"
        )
    port map (
            in0 => \N__4443\,
            in1 => \N__4465\,
            in2 => \N__4485\,
            in3 => \N__4749\,
            lcout => \fsm_ctrl_inst1.counter_dinZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5732\,
            ce => 'H',
            sr => \N__5456\
        );

    \fsm_ctrl_inst1.counter_din_1_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4746\,
            in2 => \N__4467\,
            in3 => \N__4442\,
            lcout => \fsm_ctrl_inst1.counter_dinZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5732\,
            ce => 'H',
            sr => \N__5456\
        );

    \fsm_ctrl_inst1.SEL_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4748\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \SEL_REG\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5732\,
            ce => 'H',
            sr => \N__5456\
        );

    \fsm_ctrl_inst1.SEL_RNIQ5L_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4792\,
            lcout => \fsm_ctrl_inst1.SEL_REG_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \config_register_latched_dec_inst1.DYNSR_5_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4617\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5735\,
            ce => \N__4806\,
            sr => \N__5459\
        );

    \config_register_latched_dec_inst1.DYNSR_7_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4605\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5735\,
            ce => \N__4806\,
            sr => \N__5459\
        );

    \config_register_latched_dec_inst1.DYNSR_6_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4611\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5735\,
            ce => \N__4806\,
            sr => \N__5459\
        );

    \config_register_latched_dec_inst1.STATSR_1_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4599\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5737\,
            ce => \N__5588\,
            sr => \N__5461\
        );

    \config_register_latched_dec_inst1.STATSR_2_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4593\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5737\,
            ce => \N__5588\,
            sr => \N__5461\
        );

    \config_register_latched_dec_inst1.STATSR_3_LC_6_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4587\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5738\,
            ce => \N__5587\,
            sr => \N__5462\
        );

    \config_register_latched_dec_inst1.STATSR_4_LC_6_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4581\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5738\,
            ce => \N__5587\,
            sr => \N__5462\
        );

    \config_register_latched_dec_inst1.DYNSR_12_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4821\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5733\,
            ce => \N__4815\,
            sr => \N__5457\
        );

    \config_register_latched_dec_inst1.DYNSR_13_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4869\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5733\,
            ce => \N__4815\,
            sr => \N__5457\
        );

    \config_register_latched_dec_inst1.DYNSR_15_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4851\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5733\,
            ce => \N__4815\,
            sr => \N__5457\
        );

    \config_register_latched_dec_inst1.DYNSR_14_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4857\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5733\,
            ce => \N__4815\,
            sr => \N__5457\
        );

    \config_register_latched_dec_inst1.DYNSR_9_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4839\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5736\,
            ce => \N__4814\,
            sr => \N__5460\
        );

    \config_register_latched_dec_inst1.DYNSR_8_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4845\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5736\,
            ce => \N__4814\,
            sr => \N__5460\
        );

    \config_register_latched_dec_inst1.DYNSR_10_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4833\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5736\,
            ce => \N__4814\,
            sr => \N__5460\
        );

    \config_register_latched_dec_inst1.DYNSR_11_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4827\,
            lcout => \config_register_latched_dec_inst1.DYNSRZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5736\,
            ce => \N__4814\,
            sr => \N__5460\
        );

    \config_register_latched_dec_inst1.STATSR_5_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4761\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5739\,
            ce => \N__5586\,
            sr => \N__5463\
        );

    \config_register_latched_dec_inst1.STATSR_6_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4755\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5740\,
            ce => \N__5585\,
            sr => \N__5464\
        );

    \config_register_latched_dec_inst1.STATSR_7_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4926\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5741\,
            ce => \N__5584\,
            sr => \N__5465\
        );

    \config_register_latched_dec_inst1.STATSR_8_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4920\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5741\,
            ce => \N__5584\,
            sr => \N__5465\
        );

    \config_register_latched_dec_inst1.STATSR_10_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4899\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5742\,
            ce => \N__5583\,
            sr => \N__5466\
        );

    \config_register_latched_dec_inst1.STATSR_11_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4914\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5742\,
            ce => \N__5583\,
            sr => \N__5466\
        );

    \config_register_latched_dec_inst1.STATSR_9_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4908\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5742\,
            ce => \N__5583\,
            sr => \N__5466\
        );

    \config_register_latched_dec_inst1.STATSR_13_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4887\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5744\,
            ce => \N__5582\,
            sr => \N__5468\
        );

    \config_register_latched_dec_inst1.STATSR_12_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4893\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5744\,
            ce => \N__5582\,
            sr => \N__5468\
        );

    \config_register_latched_dec_inst1.STATSR_14_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4881\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5745\,
            ce => \N__5579\,
            sr => \N__5469\
        );

    \config_register_latched_dec_inst1.STATSR_15_LC_10_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4875\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5747\,
            ce => \N__5577\,
            sr => \N__5471\
        );

    \config_register_latched_dec_inst1.STATSR_16_LC_10_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4989\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5749\,
            ce => \N__5575\,
            sr => \N__5473\
        );

    \config_register_latched_dec_inst1.STATSR_86_LC_11_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4962\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5743\,
            ce => \N__5581\,
            sr => \N__5467\
        );

    \config_register_latched_dec_inst1.STATSR_87_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4983\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5743\,
            ce => \N__5581\,
            sr => \N__5467\
        );

    \config_register_latched_dec_inst1.STATSR_85_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4956\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5743\,
            ce => \N__5581\,
            sr => \N__5467\
        );

    \config_register_latched_dec_inst1.STATSR_84_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4950\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5746\,
            ce => \N__5580\,
            sr => \N__5470\
        );

    \config_register_latched_dec_inst1.STATSR_83_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4938\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5748\,
            ce => \N__5578\,
            sr => \N__5472\
        );

    \config_register_latched_dec_inst1.STATSR_17_LC_11_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4944\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5751\,
            ce => \N__5572\,
            sr => \N__5475\
        );

    \config_register_latched_dec_inst1.STATSR_82_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4932\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5750\,
            ce => \N__5576\,
            sr => \N__5474\
        );

    \config_register_latched_dec_inst1.STATSR_81_LC_12_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5025\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5752\,
            ce => \N__5573\,
            sr => \N__5476\
        );

    \config_register_latched_dec_inst1.STATSR_18_LC_12_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5031\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5754\,
            ce => \N__5570\,
            sr => \N__5478\
        );

    \config_register_latched_dec_inst1.STATSR_80_LC_12_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5043\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5754\,
            ce => \N__5570\,
            sr => \N__5478\
        );

    \config_register_latched_dec_inst1.STATSR_34_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5019\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5753\,
            ce => \N__5574\,
            sr => \N__5477\
        );

    \config_register_latched_dec_inst1.STATSR_33_LC_13_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5013\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5753\,
            ce => \N__5574\,
            sr => \N__5477\
        );

    \config_register_latched_dec_inst1.STATSR_30_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5079\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5753\,
            ce => \N__5574\,
            sr => \N__5477\
        );

    \config_register_latched_dec_inst1.STATSR_32_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4995\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5753\,
            ce => \N__5574\,
            sr => \N__5477\
        );

    \config_register_latched_dec_inst1.STATSR_28_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5007\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5753\,
            ce => \N__5574\,
            sr => \N__5477\
        );

    \config_register_latched_dec_inst1.STATSR_27_LC_13_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5067\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5753\,
            ce => \N__5574\,
            sr => \N__5477\
        );

    \config_register_latched_dec_inst1.STATSR_31_LC_13_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5001\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5753\,
            ce => \N__5574\,
            sr => \N__5477\
        );

    \config_register_latched_dec_inst1.STATSR_29_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5085\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5753\,
            ce => \N__5574\,
            sr => \N__5477\
        );

    \config_register_latched_dec_inst1.STATSR_23_LC_13_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5139\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5755\,
            ce => \N__5571\,
            sr => \N__5479\
        );

    \config_register_latched_dec_inst1.STATSR_25_LC_13_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5049\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5755\,
            ce => \N__5571\,
            sr => \N__5479\
        );

    \config_register_latched_dec_inst1.STATSR_26_LC_13_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5073\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5755\,
            ce => \N__5571\,
            sr => \N__5479\
        );

    \config_register_latched_dec_inst1.STATSR_35_LC_13_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5061\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5755\,
            ce => \N__5571\,
            sr => \N__5479\
        );

    \config_register_latched_dec_inst1.STATSR_24_LC_13_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5055\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5755\,
            ce => \N__5571\,
            sr => \N__5479\
        );

    \config_register_latched_dec_inst1.STATSR_79_LC_13_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5151\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5756\,
            ce => \N__5568\,
            sr => \N__5480\
        );

    \config_register_latched_dec_inst1.STATSR_21_LC_13_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5127\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5756\,
            ce => \N__5568\,
            sr => \N__5480\
        );

    \config_register_latched_dec_inst1.STATSR_19_LC_13_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5037\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5756\,
            ce => \N__5568\,
            sr => \N__5480\
        );

    \config_register_latched_dec_inst1.STATSR_78_LC_13_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5109\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5756\,
            ce => \N__5568\,
            sr => \N__5480\
        );

    \config_register_latched_dec_inst1.STATSR_22_LC_13_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5145\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5756\,
            ce => \N__5568\,
            sr => \N__5480\
        );

    \config_register_latched_dec_inst1.STATSR_20_LC_13_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5133\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5756\,
            ce => \N__5568\,
            sr => \N__5480\
        );

    \config_register_latched_dec_inst1.STATSR_76_LC_13_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5121\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5758\,
            ce => \N__5566\,
            sr => \N__5482\
        );

    \config_register_latched_dec_inst1.STATSR_73_LC_13_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5211\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5758\,
            ce => \N__5566\,
            sr => \N__5482\
        );

    \config_register_latched_dec_inst1.STATSR_75_LC_13_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5097\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5758\,
            ce => \N__5566\,
            sr => \N__5482\
        );

    \config_register_latched_dec_inst1.STATSR_77_LC_13_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5115\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5758\,
            ce => \N__5566\,
            sr => \N__5482\
        );

    \config_register_latched_dec_inst1.STATSR_74_LC_13_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5103\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5758\,
            ce => \N__5566\,
            sr => \N__5482\
        );

    \config_register_latched_dec_inst1.STATSR_71_LC_13_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5181\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5760\,
            ce => \N__5564\,
            sr => \N__5484\
        );

    \config_register_latched_dec_inst1.STATSR_72_LC_13_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5091\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5760\,
            ce => \N__5564\,
            sr => \N__5484\
        );

    \config_register_latched_dec_inst1.STATSR_37_LC_14_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5199\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5757\,
            ce => \N__5569\,
            sr => \N__5481\
        );

    \config_register_latched_dec_inst1.STATSR_36_LC_14_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5205\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5757\,
            ce => \N__5569\,
            sr => \N__5481\
        );

    \config_register_latched_dec_inst1.STATSR_38_LC_14_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5193\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5757\,
            ce => \N__5569\,
            sr => \N__5481\
        );

    \config_register_latched_dec_inst1.STATSR_39_LC_14_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5187\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5757\,
            ce => \N__5569\,
            sr => \N__5481\
        );

    \config_register_latched_dec_inst1.STATSR_68_LC_14_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5169\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5762\,
            ce => \N__5561\,
            sr => \N__5486\
        );

    \config_register_latched_dec_inst1.STATSR_70_LC_14_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5157\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5762\,
            ce => \N__5561\,
            sr => \N__5486\
        );

    \config_register_latched_dec_inst1.STATSR_66_LC_14_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5277\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5762\,
            ce => \N__5561\,
            sr => \N__5486\
        );

    \config_register_latched_dec_inst1.STATSR_67_LC_14_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5175\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5762\,
            ce => \N__5561\,
            sr => \N__5486\
        );

    \config_register_latched_dec_inst1.STATSR_69_LC_14_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5163\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5762\,
            ce => \N__5561\,
            sr => \N__5486\
        );

    \config_register_latched_dec_inst1.STATSR_40_LC_15_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5253\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5759\,
            ce => \N__5567\,
            sr => \N__5483\
        );

    \config_register_latched_dec_inst1.STATSR_41_LC_15_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5247\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5759\,
            ce => \N__5567\,
            sr => \N__5483\
        );

    \config_register_latched_dec_inst1.STATSR_43_LC_15_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5235\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5759\,
            ce => \N__5567\,
            sr => \N__5483\
        );

    \config_register_latched_dec_inst1.STATSR_42_LC_15_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5241\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5759\,
            ce => \N__5567\,
            sr => \N__5483\
        );

    \config_register_latched_dec_inst1.STATSR_44_LC_15_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5229\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5759\,
            ce => \N__5567\,
            sr => \N__5483\
        );

    \config_register_latched_dec_inst1.STATSR_57_LC_15_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5784\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5763\,
            ce => \N__5562\,
            sr => \N__5487\
        );

    \config_register_latched_dec_inst1.STATSR_61_LC_15_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5217\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5763\,
            ce => \N__5562\,
            sr => \N__5487\
        );

    \config_register_latched_dec_inst1.STATSR_59_LC_15_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5307\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5763\,
            ce => \N__5562\,
            sr => \N__5487\
        );

    \config_register_latched_dec_inst1.STATSR_60_LC_15_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5223\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5763\,
            ce => \N__5562\,
            sr => \N__5487\
        );

    \config_register_latched_dec_inst1.STATSR_58_LC_15_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5313\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5763\,
            ce => \N__5562\,
            sr => \N__5487\
        );

    \config_register_latched_dec_inst1.STATSR_64_LC_15_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5289\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5765\,
            ce => \N__5559\,
            sr => \N__5489\
        );

    \config_register_latched_dec_inst1.STATSR_62_LC_15_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5301\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5765\,
            ce => \N__5559\,
            sr => \N__5489\
        );

    \config_register_latched_dec_inst1.STATSR_63_LC_15_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5295\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5765\,
            ce => \N__5559\,
            sr => \N__5489\
        );

    \config_register_latched_dec_inst1.STATSR_65_LC_15_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5283\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5765\,
            ce => \N__5559\,
            sr => \N__5489\
        );

    \config_register_latched_dec_inst1.STATSR_47_LC_16_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5271\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5761\,
            ce => \N__5565\,
            sr => \N__5485\
        );

    \config_register_latched_dec_inst1.STATSR_46_LC_16_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5259\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5761\,
            ce => \N__5565\,
            sr => \N__5485\
        );

    \config_register_latched_dec_inst1.STATSR_45_LC_16_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5265\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5761\,
            ce => \N__5565\,
            sr => \N__5485\
        );

    \config_register_latched_dec_inst1.STATSR_51_LC_16_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5808\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5764\,
            ce => \N__5563\,
            sr => \N__5488\
        );

    \config_register_latched_dec_inst1.STATSR_48_LC_16_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5826\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5764\,
            ce => \N__5563\,
            sr => \N__5488\
        );

    \config_register_latched_dec_inst1.STATSR_49_LC_16_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5820\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5764\,
            ce => \N__5563\,
            sr => \N__5488\
        );

    \config_register_latched_dec_inst1.STATSR_50_LC_16_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5814\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5764\,
            ce => \N__5563\,
            sr => \N__5488\
        );

    \config_register_latched_dec_inst1.STATSR_52_LC_16_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5802\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5764\,
            ce => \N__5563\,
            sr => \N__5488\
        );

    \config_register_latched_dec_inst1.STATSR_54_LC_16_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5790\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5764\,
            ce => \N__5563\,
            sr => \N__5488\
        );

    \config_register_latched_dec_inst1.STATSR_53_LC_16_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5796\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5764\,
            ce => \N__5563\,
            sr => \N__5488\
        );

    \config_register_latched_dec_inst1.STATSR_56_LC_16_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5772\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5766\,
            ce => \N__5560\,
            sr => \N__5490\
        );

    \config_register_latched_dec_inst1.STATSR_55_LC_16_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5778\,
            lcout => \config_register_latched_dec_inst1.STATSRZ0Z_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5766\,
            ce => \N__5560\,
            sr => \N__5490\
        );
end \INTERFACE\;
